
module controller ( clk, rst_n, test_mode, operation, apnpsf_complete, 
        apnpsf_en, complete );
  input [2:0] operation;
  input clk, rst_n, test_mode, apnpsf_complete;
  output apnpsf_en, complete;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [1:0] state;
  wire   [1:0] next_state;

  DFFARX1 next_state_reg_0_ ( .D(n14), .CLK(clk), .RSTB(rst_n), .Q(
        next_state[0]), .QN(n4) );
  DFFASX1 state_reg_0_ ( .D(n4), .CLK(clk), .SETB(rst_n), .QN(state[0]) );
  DFFARX1 next_state_reg_1_ ( .D(n13), .CLK(clk), .RSTB(rst_n), .Q(
        next_state[1]), .QN(n2) );
  DFFASX1 state_reg_1_ ( .D(n2), .CLK(clk), .SETB(rst_n), .Q(n5), .QN(state[1]) );
  DFFARX1 apnpsf_en_reg ( .D(n12), .CLK(clk), .RSTB(rst_n), .Q(apnpsf_en) );
  OA21X1 U3 ( .IN1(state[0]), .IN2(apnpsf_en), .IN3(state[1]), .Q(n12) );
  NAND3X0 U6 ( .IN1(n9), .IN2(n10), .IN3(n7), .QN(n14) );
  NOR2X0 U10 ( .IN1(state[0]), .IN2(n5), .QN(n8) );
  NAND2X0 U8 ( .IN1(apnpsf_complete), .IN2(state[1]), .QN(n11) );
  NAND2X0 U7 ( .IN1(n11), .IN2(state[0]), .QN(n7) );
  NAND2X0 U11 ( .IN1(n5), .IN2(test_mode), .QN(n9) );
  NAND2X0 U9 ( .IN1(n8), .IN2(next_state[0]), .QN(n10) );
  NAND2X0 U5 ( .IN1(n8), .IN2(next_state[1]), .QN(n6) );
  NAND2X0 U4 ( .IN1(n6), .IN2(n7), .QN(n13) );
  NBUFFX2 U12 ( .IN(apnpsf_complete), .Q(complete) );
endmodule


module apnpsf_controller ( clk, rst_n, apnpsf_en, memtype, address, counter, 
        start, en1, en2, en3, en4, en5, en6, en7, en8, en9, en10, en11, en12, 
        en13, en14, en15, en16, finish );
  input [4:0] memtype;
  input [15:0] address;
  input [8:0] counter;
  input clk, rst_n, apnpsf_en;
  output start, en1, en2, en3, en4, en5, en6, en7, en8, en9, en10, en11, en12,
         en13, en14, en15, en16, finish;
  wire   n18, n19, n20, n22, n23, n35, n36, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n21, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130;
  wire   [4:0] apnpsf_state;
  wire   [4:0] next_apnpsf;

  DFFARX1 finish_reg ( .D(n182), .CLK(clk), .RSTB(rst_n), .Q(finish) );
  DFFARX1 next_apnpsf_reg_1_ ( .D(n180), .CLK(clk), .RSTB(rst_n), .Q(
        next_apnpsf[1]), .QN(n23) );
  DFFASX1 apnpsf_state_reg_1_ ( .D(n23), .CLK(clk), .SETB(rst_n), .Q(n21), 
        .QN(apnpsf_state[1]) );
  DFFARX1 next_apnpsf_reg_0_ ( .D(n181), .CLK(clk), .RSTB(rst_n), .Q(
        next_apnpsf[0]), .QN(n22) );
  DFFARX1 next_apnpsf_reg_2_ ( .D(n179), .CLK(clk), .RSTB(rst_n), .Q(
        next_apnpsf[2]), .QN(n20) );
  DFFASX1 apnpsf_state_reg_2_ ( .D(n20), .CLK(clk), .SETB(rst_n), .Q(n36), 
        .QN(n25) );
  DFFARX1 next_apnpsf_reg_4_ ( .D(n178), .CLK(clk), .RSTB(rst_n), .Q(
        next_apnpsf[4]), .QN(n19) );
  DFFASX1 apnpsf_state_reg_4_ ( .D(n19), .CLK(clk), .SETB(rst_n), .Q(n26), 
        .QN(apnpsf_state[4]) );
  DFFARX1 next_apnpsf_reg_3_ ( .D(n177), .CLK(clk), .RSTB(rst_n), .Q(
        next_apnpsf[3]), .QN(n18) );
  DFFASX1 apnpsf_state_reg_3_ ( .D(n18), .CLK(clk), .SETB(rst_n), .Q(n35), 
        .QN(n27) );
  DFFARX1 en16_reg ( .D(n175), .CLK(clk), .RSTB(rst_n), .Q(en16) );
  DFFARX1 start_reg ( .D(n176), .CLK(clk), .RSTB(rst_n), .Q(start) );
  DFFARX1 en1_reg ( .D(n174), .CLK(clk), .RSTB(rst_n), .Q(en1) );
  DFFARX1 en2_reg ( .D(n173), .CLK(clk), .RSTB(rst_n), .Q(en2) );
  DFFARX1 en3_reg ( .D(n172), .CLK(clk), .RSTB(rst_n), .Q(en3) );
  DFFARX1 en4_reg ( .D(n171), .CLK(clk), .RSTB(rst_n), .Q(en4) );
  DFFARX1 en5_reg ( .D(n170), .CLK(clk), .RSTB(rst_n), .Q(en5) );
  DFFARX1 en6_reg ( .D(n169), .CLK(clk), .RSTB(rst_n), .Q(en6) );
  DFFARX1 en7_reg ( .D(n168), .CLK(clk), .RSTB(rst_n), .Q(en7) );
  DFFARX1 en8_reg ( .D(n167), .CLK(clk), .RSTB(rst_n), .Q(en8) );
  DFFARX1 en9_reg ( .D(n166), .CLK(clk), .RSTB(rst_n), .Q(en9) );
  DFFARX1 en10_reg ( .D(n165), .CLK(clk), .RSTB(rst_n), .Q(en10) );
  DFFARX1 en11_reg ( .D(n164), .CLK(clk), .RSTB(rst_n), .Q(en11) );
  DFFARX1 en12_reg ( .D(n163), .CLK(clk), .RSTB(rst_n), .Q(en12) );
  DFFARX1 en13_reg ( .D(n162), .CLK(clk), .RSTB(rst_n), .Q(en13) );
  DFFARX1 en14_reg ( .D(n161), .CLK(clk), .RSTB(rst_n), .Q(en14) );
  DFFARX1 en15_reg ( .D(n160), .CLK(clk), .RSTB(rst_n), .Q(en15) );
  DFFASX1 apnpsf_state_reg_0_ ( .D(n22), .CLK(clk), .SETB(rst_n), .Q(n28), 
        .QN(apnpsf_state[0]) );
  NAND2X0 U3 ( .IN1(n119), .IN2(n91), .QN(n85) );
  NAND2X0 U4 ( .IN1(n71), .IN2(n52), .QN(n68) );
  NAND2X0 U5 ( .IN1(n113), .IN2(n104), .QN(n73) );
  NAND2X0 U6 ( .IN1(n65), .IN2(n64), .QN(n76) );
  NAND2X0 U7 ( .IN1(n65), .IN2(n57), .QN(n104) );
  NAND2X0 U8 ( .IN1(n58), .IN2(n57), .QN(n51) );
  NAND2X0 U9 ( .IN1(next_apnpsf[3]), .IN2(n102), .QN(n103) );
  NAND2X0 U10 ( .IN1(next_apnpsf[4]), .IN2(n102), .QN(n97) );
  NAND2X0 U11 ( .IN1(n119), .IN2(n123), .QN(n77) );
  NAND2X0 U12 ( .IN1(n130), .IN2(n129), .QN(n160) );
  NAND2X0 U13 ( .IN1(n127), .IN2(n126), .QN(n161) );
  NAND2X0 U14 ( .IN1(n118), .IN2(n117), .QN(n167) );
  NAND2X0 U15 ( .IN1(n116), .IN2(n115), .QN(n168) );
  NAND2X0 U16 ( .IN1(n110), .IN2(n109), .QN(n175) );
  NAND2X0 U17 ( .IN1(en8), .IN2(n128), .QN(n118) );
  NAND2X0 U18 ( .IN1(en14), .IN2(n128), .QN(n127) );
  NAND2X0 U19 ( .IN1(en15), .IN2(n128), .QN(n130) );
  NAND2X0 U20 ( .IN1(n120), .IN2(n123), .QN(n126) );
  NAND2X0 U21 ( .IN1(n124), .IN2(n121), .QN(n117) );
  NAND3X0 U22 ( .IN1(n124), .IN2(n112), .IN3(apnpsf_en), .QN(n83) );
  NAND2X0 U23 ( .IN1(n36), .IN2(n35), .QN(n55) );
  NAND2X0 U24 ( .IN1(n21), .IN2(n26), .QN(n86) );
  OA221X1 U25 ( .IN1(n55), .IN2(apnpsf_state[1]), .IN3(n55), .IN4(
        apnpsf_state[0]), .IN5(apnpsf_state[4]), .Q(n128) );
  NAND2X0 U26 ( .IN1(n35), .IN2(n90), .QN(n115) );
  NAND2X0 U27 ( .IN1(n90), .IN2(n27), .QN(n129) );
  NOR2X0 U28 ( .IN1(n35), .IN2(n25), .QN(n121) );
  NOR2X0 U29 ( .IN1(apnpsf_state[0]), .IN2(n86), .QN(n124) );
  NOR2X0 U30 ( .IN1(n25), .IN2(n27), .QN(n112) );
  NAND2X0 U31 ( .IN1(n35), .IN2(n25), .QN(n88) );
  NAND2X0 U32 ( .IN1(n25), .IN2(n27), .QN(n87) );
  NOR2X0 U33 ( .IN1(apnpsf_state[0]), .IN2(n56), .QN(n120) );
  NAND2X0 U34 ( .IN1(apnpsf_state[1]), .IN2(n26), .QN(n56) );
  INVX0 U35 ( .IN(n69), .QN(n119) );
  NAND2X0 U36 ( .IN1(apnpsf_state[0]), .IN2(n89), .QN(n69) );
  AO22X1 U37 ( .IN1(n120), .IN2(n112), .IN3(en2), .IN4(n128), .Q(n173) );
  AO22X1 U38 ( .IN1(n119), .IN2(n121), .IN3(en9), .IN4(n128), .Q(n166) );
  AO22X1 U39 ( .IN1(n124), .IN2(n123), .IN3(en12), .IN4(n128), .Q(n163) );
  AO22X1 U40 ( .IN1(n119), .IN2(n112), .IN3(en1), .IN4(n128), .Q(n174) );
  AO22X1 U41 ( .IN1(n122), .IN2(n112), .IN3(en3), .IN4(n128), .Q(n172) );
  AO22X1 U42 ( .IN1(n114), .IN2(n124), .IN3(en4), .IN4(n128), .Q(n171) );
  AO22X1 U43 ( .IN1(n114), .IN2(n120), .IN3(en6), .IN4(n128), .Q(n169) );
  AO22X1 U44 ( .IN1(n122), .IN2(n121), .IN3(en11), .IN4(n128), .Q(n164) );
  AO22X1 U45 ( .IN1(n120), .IN2(n121), .IN3(en10), .IN4(n128), .Q(n165) );
  NAND4X0 U46 ( .IN1(apnpsf_state[4]), .IN2(apnpsf_state[0]), .IN3(n112), 
        .IN4(n21), .QN(n54) );
  INVX0 U47 ( .IN(n54), .QN(n62) );
  AO21X1 U48 ( .IN1(finish), .IN2(n128), .IN3(n62), .Q(n182) );
  INVX0 U49 ( .IN(address[1]), .QN(n52) );
  AND3X1 U50 ( .IN1(counter[0]), .IN2(counter[3]), .IN3(counter[1]), .Q(n29)
         );
  AND3X1 U51 ( .IN1(counter[2]), .IN2(counter[4]), .IN3(n29), .Q(n30) );
  OR3X1 U52 ( .IN1(n30), .IN2(counter[6]), .IN3(counter[5]), .Q(n31) );
  AND3X1 U53 ( .IN1(counter[8]), .IN2(counter[7]), .IN3(n31), .Q(n58) );
  AND3X1 U54 ( .IN1(n52), .IN2(address[0]), .IN3(n58), .Q(n65) );
  AND4X1 U55 ( .IN1(address[4]), .IN2(address[6]), .IN3(address[8]), .IN4(
        address[7]), .Q(n32) );
  NAND4X0 U56 ( .IN1(address[5]), .IN2(address[2]), .IN3(address[3]), .IN4(n32), .QN(n40) );
  INVX0 U57 ( .IN(n40), .QN(n33) );
  NAND3X0 U58 ( .IN1(n33), .IN2(address[10]), .IN3(address[9]), .QN(n38) );
  INVX0 U59 ( .IN(n38), .QN(n34) );
  NAND3X0 U60 ( .IN1(n34), .IN2(address[11]), .IN3(address[12]), .QN(n43) );
  INVX0 U61 ( .IN(n43), .QN(n37) );
  NAND3X0 U62 ( .IN1(n37), .IN2(address[13]), .IN3(address[14]), .QN(n50) );
  INVX0 U63 ( .IN(memtype[2]), .QN(n42) );
  NOR2X0 U64 ( .IN1(address[11]), .IN2(n42), .QN(n39) );
  NOR3X0 U65 ( .IN1(n39), .IN2(memtype[4]), .IN3(n38), .QN(n49) );
  NOR2X0 U66 ( .IN1(address[9]), .IN2(n42), .QN(n41) );
  NOR4X0 U67 ( .IN1(n41), .IN2(memtype[4]), .IN3(memtype[3]), .IN4(n40), .QN(
        n48) );
  NOR2X0 U68 ( .IN1(address[13]), .IN2(n42), .QN(n44) );
  NOR3X0 U69 ( .IN1(n44), .IN2(memtype[3]), .IN3(n43), .QN(n47) );
  INVX0 U70 ( .IN(address[15]), .QN(n45) );
  NOR2X0 U71 ( .IN1(n50), .IN2(n45), .QN(n46) );
  NOR4X0 U72 ( .IN1(n49), .IN2(n48), .IN3(n47), .IN4(n46), .QN(n63) );
  OAI21X1 U73 ( .IN1(memtype[2]), .IN2(n50), .IN3(n63), .QN(n57) );
  NOR2X0 U74 ( .IN1(n36), .IN2(n104), .QN(n53) );
  NOR2X0 U75 ( .IN1(address[0]), .IN2(n51), .QN(n71) );
  NOR2X0 U76 ( .IN1(n25), .IN2(n68), .QN(n91) );
  NAND3X0 U77 ( .IN1(apnpsf_state[1]), .IN2(apnpsf_state[0]), .IN3(n26), .QN(
        n111) );
  NOR3X0 U78 ( .IN1(n53), .IN2(n91), .IN3(n111), .QN(n80) );
  NOR2X0 U79 ( .IN1(finish), .IN2(n54), .QN(n98) );
  NOR4X0 U80 ( .IN1(apnpsf_state[0]), .IN2(n26), .IN3(n21), .IN4(n55), .QN(
        n108) );
  NAND4X0 U81 ( .IN1(apnpsf_state[4]), .IN2(n112), .IN3(n21), .IN4(n28), .QN(
        n109) );
  NAND2X0 U82 ( .IN1(n120), .IN2(n25), .QN(n94) );
  NAND3X0 U83 ( .IN1(n117), .IN2(n109), .IN3(n94), .QN(n61) );
  AND3X1 U84 ( .IN1(address[0]), .IN2(address[1]), .IN3(n57), .Q(n82) );
  OA221X1 U85 ( .IN1(n108), .IN2(n58), .IN3(n108), .IN4(n61), .IN5(n82), .Q(
        n67) );
  NOR3X0 U86 ( .IN1(n36), .IN2(n21), .IN3(apnpsf_state[0]), .QN(n59) );
  NOR2X0 U87 ( .IN1(n59), .IN2(apnpsf_state[4]), .QN(n60) );
  NOR4X0 U88 ( .IN1(n62), .IN2(n108), .IN3(n61), .IN4(n60), .QN(n102) );
  INVX0 U89 ( .IN(n86), .QN(n89) );
  INVX0 U90 ( .IN(n87), .QN(n123) );
  INVX0 U91 ( .IN(n77), .QN(n125) );
  INVX0 U92 ( .IN(n63), .QN(n64) );
  AO22X1 U93 ( .IN1(n102), .IN2(next_apnpsf[0]), .IN3(n125), .IN4(n76), .Q(n66) );
  NOR4X0 U94 ( .IN1(n80), .IN2(n98), .IN3(n67), .IN4(n66), .QN(n75) );
  NAND3X0 U95 ( .IN1(n36), .IN2(n119), .IN3(n68), .QN(n74) );
  NOR2X0 U96 ( .IN1(n69), .IN2(n88), .QN(n113) );
  MUX21X1 U97 ( .IN1(n124), .IN2(n120), .S(n36), .Q(n70) );
  NAND3X0 U98 ( .IN1(n71), .IN2(address[1]), .IN3(n70), .QN(n72) );
  NAND4X0 U99 ( .IN1(n75), .IN2(n74), .IN3(n73), .IN4(n72), .QN(n181) );
  NOR2X0 U100 ( .IN1(n77), .IN2(n76), .QN(n79) );
  INVX0 U101 ( .IN(n104), .QN(n93) );
  AO22X1 U102 ( .IN1(n93), .IN2(n113), .IN3(n102), .IN4(next_apnpsf[1]), .Q(
        n78) );
  NOR4X0 U103 ( .IN1(n80), .IN2(n120), .IN3(n79), .IN4(n78), .QN(n84) );
  INVX0 U104 ( .IN(n108), .QN(n81) );
  OA22X1 U105 ( .IN1(finish), .IN2(n83), .IN3(n82), .IN4(n81), .Q(n101) );
  NAND3X0 U106 ( .IN1(n85), .IN2(n84), .IN3(n101), .QN(n180) );
  NOR2X0 U107 ( .IN1(n36), .IN2(n111), .QN(n90) );
  OA22X1 U108 ( .IN1(n93), .IN2(n129), .IN3(n87), .IN4(n86), .Q(n107) );
  INVX0 U109 ( .IN(n88), .QN(n114) );
  AOI22X1 U110 ( .IN1(n89), .IN2(n114), .IN3(n102), .IN4(next_apnpsf[2]), .QN(
        n96) );
  INVX0 U111 ( .IN(n91), .QN(n92) );
  OA22X1 U112 ( .IN1(n93), .IN2(n115), .IN3(n111), .IN4(n92), .Q(n95) );
  NAND4X0 U113 ( .IN1(n107), .IN2(n96), .IN3(n95), .IN4(n94), .QN(n179) );
  OA21X1 U114 ( .IN1(n129), .IN2(n104), .IN3(n97), .Q(n100) );
  INVX0 U115 ( .IN(n98), .QN(n99) );
  NAND4X0 U116 ( .IN1(n101), .IN2(n100), .IN3(n99), .IN4(n109), .QN(n178) );
  OA21X1 U117 ( .IN1(n115), .IN2(n104), .IN3(n103), .Q(n106) );
  NAND2X0 U118 ( .IN1(n121), .IN2(n26), .QN(n105) );
  NAND4X0 U119 ( .IN1(n107), .IN2(n106), .IN3(n105), .IN4(n126), .QN(n177) );
  AO21X1 U120 ( .IN1(start), .IN2(n128), .IN3(n108), .Q(n176) );
  NAND2X0 U121 ( .IN1(en16), .IN2(n128), .QN(n110) );
  INVX0 U122 ( .IN(n111), .QN(n122) );
  AO21X1 U123 ( .IN1(en5), .IN2(n128), .IN3(n113), .Q(n170) );
  NAND2X0 U124 ( .IN1(en7), .IN2(n128), .QN(n116) );
  AO21X1 U125 ( .IN1(en13), .IN2(n128), .IN3(n125), .Q(n162) );
endmodule


module apnpsf_datapath ( clk, rst_n, start, en1, en2, en3, en4, en5, en6, en7, 
        en8, en9, en10, en11, en12, en13, en14, en15, en16, 
        error_exceed_ignore, allowable_faulty, address, write_read, wdata, 
        rdata, counter, error, force_terminate, memtype );
  input [15:0] allowable_faulty;
  output [15:0] address;
  output [63:0] wdata;
  input [63:0] rdata;
  output [8:0] counter;
  input [4:0] memtype;
  input clk, rst_n, start, en1, en2, en3, en4, en5, en6, en7, en8, en9, en10,
         en11, en12, en13, en14, en15, en16, error_exceed_ignore;
  output write_read, error, force_terminate;
  wire   N111, N112, N113, N114, N115, N116, N117, N118, N119, N133, N134,
         N135, N136, N137, N138, N139, N140, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, write_read_2, N255, N256,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, C36_DATA3_0, C36_DATA3_1, C36_DATA3_2, C36_DATA3_3,
         C36_DATA3_4, C36_DATA3_5, C36_DATA3_6, C36_DATA3_7, C36_DATA3_8,
         C36_DATA3_9, C36_DATA3_10, C36_DATA3_11, C36_DATA3_12, C36_DATA3_13,
         C36_DATA3_14, n203, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851,
         RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_2,
         RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_1,
         DP_OP_350_296_6706_n40, DP_OP_350_296_6706_n22,
         DP_OP_350_296_6706_n21, DP_OP_350_296_6706_n16,
         DP_OP_350_296_6706_n15, DP_OP_350_296_6706_n14,
         DP_OP_350_296_6706_n13, DP_OP_350_296_6706_n12,
         DP_OP_350_296_6706_n11, DP_OP_350_296_6706_n10, DP_OP_350_296_6706_n9,
         DP_OP_350_296_6706_n8, DP_OP_350_296_6706_n7, DP_OP_350_296_6706_n6,
         DP_OP_350_296_6706_n5, DP_OP_350_296_6706_n4, DP_OP_350_296_6706_n3,
         DP_OP_350_296_6706_n2, n1, n2, n3, n4, n5, n6, n7, n8, n9, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n100, n102, n104, n106, n107, n109, n111, n112, n113, n116, n117,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917;
  wire   [7:0] counter_1;
  wire   [63:0] wdata_2;
  wire   [63:0] rdata_cp;
  wire   [15:0] address_1;
  wire   [15:0] address_2;
  wire   [15:0] error_counter;

  DFFARX1 counter_reg_0_ ( .D(N111), .CLK(clk), .RSTB(rst_n), .Q(counter[0]), 
        .QN(n244) );
  DFFARX1 counter_reg_8_ ( .D(N119), .CLK(clk), .RSTB(rst_n), .Q(counter[8]), 
        .QN(n238) );
  DFFARX1 counter_reg_7_ ( .D(N118), .CLK(clk), .RSTB(rst_n), .Q(counter[7]), 
        .QN(n232) );
  DFFARX1 counter_reg_6_ ( .D(N117), .CLK(clk), .RSTB(rst_n), .Q(counter[6]), 
        .QN(n234) );
  DFFARX1 counter_reg_5_ ( .D(N116), .CLK(clk), .RSTB(rst_n), .Q(counter[5]), 
        .QN(n237) );
  DFFARX1 counter_reg_4_ ( .D(N115), .CLK(clk), .RSTB(rst_n), .Q(counter[4]), 
        .QN(n235) );
  DFFARX1 counter_reg_3_ ( .D(N114), .CLK(clk), .RSTB(rst_n), .Q(counter[3]), 
        .QN(n245) );
  DFFARX1 counter_reg_2_ ( .D(N113), .CLK(clk), .RSTB(rst_n), .Q(counter[2]), 
        .QN(n236) );
  DFFARX1 counter_reg_1_ ( .D(N112), .CLK(clk), .RSTB(rst_n), .Q(counter[1]), 
        .QN(n233) );
  DFFARX1 rdata_cp_reg_7_ ( .D(rdata[7]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[7]) );
  DFFARX1 rdata_cp_reg_6_ ( .D(rdata[6]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[6]) );
  DFFARX1 rdata_cp_reg_5_ ( .D(rdata[5]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[5]) );
  DFFARX1 rdata_cp_reg_4_ ( .D(rdata[4]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[4]) );
  DFFARX1 rdata_cp_reg_3_ ( .D(rdata[3]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[3]) );
  DFFARX1 rdata_cp_reg_2_ ( .D(rdata[2]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[2]) );
  DFFARX1 rdata_cp_reg_1_ ( .D(rdata[1]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[1]) );
  DFFARX1 rdata_cp_reg_0_ ( .D(rdata[0]), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[0]) );
  DFFARX1 counter_1_reg_7_ ( .D(N140), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[7]), .QN(n337) );
  DFFARX1 counter_1_reg_6_ ( .D(N139), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[6]), .QN(n328) );
  DFFARX1 counter_1_reg_5_ ( .D(N138), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[5]) );
  DFFARX1 counter_1_reg_4_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[4]), .QN(n327) );
  DFFARX1 counter_1_reg_3_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[3]), .QN(n255) );
  DFFARX1 counter_1_reg_2_ ( .D(N135), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[2]), .QN(n260) );
  DFFARX1 counter_1_reg_1_ ( .D(N134), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[1]) );
  DFFARX1 counter_1_reg_0_ ( .D(N133), .CLK(clk), .RSTB(rst_n), .Q(
        counter_1[0]) );
  DFFARX1 address_1_reg_0_ ( .D(N255), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[0]), .QN(n261) );
  DFFARX1 address_1_reg_15_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[15]), .QN(n333) );
  DFFARX1 address_1_reg_14_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[14]) );
  DFFARX1 address_1_reg_13_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[13]), .QN(n247) );
  DFFARX1 address_1_reg_12_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[12]) );
  DFFARX1 address_1_reg_11_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[11]), .QN(n259) );
  DFFARX1 address_1_reg_10_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[10]) );
  DFFARX1 address_1_reg_9_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[9]), .QN(n262) );
  DFFARX1 address_1_reg_8_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[8]), .QN(n250) );
  DFFARX1 address_1_reg_7_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[7]) );
  DFFARX1 address_1_reg_6_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[6]), .QN(n249) );
  DFFARX1 address_1_reg_5_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[5]) );
  DFFARX1 address_1_reg_4_ ( .D(N259), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[4]), .QN(n252) );
  DFFARX1 address_1_reg_3_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[3]) );
  DFFARX1 address_1_reg_2_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[2]), .QN(n336) );
  DFFARX1 address_1_reg_1_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[1]) );
  DFFARX1 error_counter_reg_15_ ( .D(n754), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[15]), .QN(n241) );
  DFFARX1 error_counter_reg_14_ ( .D(n755), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[14]), .QN(n335) );
  DFFARX1 error_counter_reg_13_ ( .D(n756), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[13]), .QN(n257) );
  DFFARX1 error_counter_reg_12_ ( .D(n757), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[12]), .QN(n334) );
  DFFARX1 error_counter_reg_11_ ( .D(n758), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[11]), .QN(n240) );
  DFFARX1 error_counter_reg_10_ ( .D(n759), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[10]), .QN(n332) );
  DFFARX1 error_counter_reg_9_ ( .D(n760), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[9]), .QN(n242) );
  DFFARX1 error_counter_reg_8_ ( .D(n761), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[8]), .QN(n329) );
  DFFARX1 error_counter_reg_7_ ( .D(n762), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[7]), .QN(n243) );
  DFFARX1 error_counter_reg_6_ ( .D(n763), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[6]), .QN(n331) );
  DFFARX1 error_counter_reg_5_ ( .D(n764), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[5]), .QN(n258) );
  DFFARX1 error_counter_reg_4_ ( .D(n765), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[4]), .QN(n330) );
  DFFARX1 error_counter_reg_3_ ( .D(n766), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[3]), .QN(n248) );
  DFFARX1 error_counter_reg_2_ ( .D(n767), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[2]), .QN(n253) );
  DFFARX1 error_counter_reg_1_ ( .D(n768), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[1]), .QN(n239) );
  DFFARX1 error_counter_reg_0_ ( .D(n769), .CLK(clk), .RSTB(rst_n), .Q(
        error_counter[0]), .QN(n251) );
  DFFARX1 write_read_2_reg ( .D(n851), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_2) );
  DFFARX1 address_2_reg_0_ ( .D(n850), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[0]) );
  DFFARX1 address_2_reg_1_ ( .D(n849), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[1]) );
  DFFARX1 address_2_reg_2_ ( .D(n848), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[2]) );
  DFFARX1 address_2_reg_3_ ( .D(n847), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[3]) );
  DFFARX1 address_2_reg_4_ ( .D(n846), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[4]) );
  DFFARX1 address_2_reg_5_ ( .D(n845), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[5]) );
  DFFARX1 address_2_reg_6_ ( .D(n844), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[6]) );
  DFFARX1 address_2_reg_7_ ( .D(n843), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[7]) );
  DFFARX1 address_2_reg_8_ ( .D(n842), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[8]) );
  DFFARX1 address_2_reg_9_ ( .D(n841), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[9]) );
  DFFARX1 address_2_reg_10_ ( .D(n840), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[10]) );
  DFFARX1 address_2_reg_11_ ( .D(n839), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[11]) );
  DFFARX1 address_2_reg_12_ ( .D(n838), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[12]) );
  DFFARX1 address_2_reg_13_ ( .D(n837), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[13]) );
  DFFARX1 address_2_reg_14_ ( .D(n836), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[14]) );
  DFFARX1 address_2_reg_15_ ( .D(n835), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[15]) );
  DFFARX1 wdata_2_reg_63_ ( .D(n834), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[63]), 
        .QN(n300) );
  DFFARX1 rdata_cp_reg_63_ ( .D(N200), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[63]) );
  DFFARX1 wdata_2_reg_62_ ( .D(n833), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[62]), 
        .QN(n263) );
  DFFARX1 rdata_cp_reg_62_ ( .D(N199), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[62]) );
  DFFARX1 wdata_2_reg_61_ ( .D(n832), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[61]), 
        .QN(n299) );
  DFFARX1 rdata_cp_reg_61_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[61]) );
  DFFARX1 wdata_2_reg_60_ ( .D(n831), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[60]), 
        .QN(n298) );
  DFFARX1 rdata_cp_reg_60_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[60]) );
  DFFARX1 wdata_2_reg_59_ ( .D(n830), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[59]), 
        .QN(n297) );
  DFFARX1 rdata_cp_reg_59_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[59]) );
  DFFARX1 wdata_2_reg_58_ ( .D(n829), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[58]), 
        .QN(n296) );
  DFFARX1 rdata_cp_reg_58_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[58]) );
  DFFARX1 wdata_2_reg_57_ ( .D(n828), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[57]), 
        .QN(n295) );
  DFFARX1 rdata_cp_reg_57_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[57]) );
  DFFARX1 wdata_2_reg_56_ ( .D(n827), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[56]), 
        .QN(n294) );
  DFFARX1 rdata_cp_reg_56_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[56]) );
  DFFARX1 wdata_2_reg_55_ ( .D(n826), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[55]), 
        .QN(n293) );
  DFFARX1 rdata_cp_reg_55_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[55]) );
  DFFARX1 wdata_2_reg_54_ ( .D(n825), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[54]), 
        .QN(n292) );
  DFFARX1 rdata_cp_reg_54_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[54]) );
  DFFARX1 wdata_2_reg_53_ ( .D(n824), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[53]), 
        .QN(n291) );
  DFFARX1 rdata_cp_reg_53_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[53]) );
  DFFARX1 wdata_2_reg_52_ ( .D(n823), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[52]), 
        .QN(n290) );
  DFFARX1 rdata_cp_reg_52_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[52]) );
  DFFARX1 wdata_2_reg_51_ ( .D(n822), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[51]), 
        .QN(n289) );
  DFFARX1 rdata_cp_reg_51_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[51]) );
  DFFARX1 wdata_2_reg_50_ ( .D(n821), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[50]), 
        .QN(n288) );
  DFFARX1 rdata_cp_reg_50_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[50]) );
  DFFARX1 wdata_2_reg_49_ ( .D(n820), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[49]), 
        .QN(n287) );
  DFFARX1 rdata_cp_reg_49_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[49]) );
  DFFARX1 wdata_2_reg_48_ ( .D(n819), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[48]), 
        .QN(n286) );
  DFFARX1 rdata_cp_reg_48_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[48]) );
  DFFARX1 wdata_2_reg_47_ ( .D(n818), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[47]), 
        .QN(n285) );
  DFFARX1 rdata_cp_reg_47_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[47]) );
  DFFARX1 wdata_2_reg_46_ ( .D(n817), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[46]), 
        .QN(n284) );
  DFFARX1 rdata_cp_reg_46_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[46]) );
  DFFARX1 wdata_2_reg_45_ ( .D(n816), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[45]), 
        .QN(n283) );
  DFFARX1 rdata_cp_reg_45_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[45]) );
  DFFARX1 wdata_2_reg_44_ ( .D(n815), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[44]), 
        .QN(n282) );
  DFFARX1 rdata_cp_reg_44_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[44]) );
  DFFARX1 wdata_2_reg_43_ ( .D(n814), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[43]), 
        .QN(n281) );
  DFFARX1 rdata_cp_reg_43_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[43]) );
  DFFARX1 wdata_2_reg_42_ ( .D(n813), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[42]), 
        .QN(n280) );
  DFFARX1 rdata_cp_reg_42_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[42]) );
  DFFARX1 wdata_2_reg_41_ ( .D(n812), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[41]), 
        .QN(n279) );
  DFFARX1 rdata_cp_reg_41_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[41]) );
  DFFARX1 wdata_2_reg_40_ ( .D(n811), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[40]), 
        .QN(n278) );
  DFFARX1 rdata_cp_reg_40_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[40]) );
  DFFARX1 wdata_2_reg_39_ ( .D(n810), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[39]), 
        .QN(n277) );
  DFFARX1 rdata_cp_reg_39_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[39]) );
  DFFARX1 wdata_2_reg_38_ ( .D(n809), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[38]), 
        .QN(n276) );
  DFFARX1 rdata_cp_reg_38_ ( .D(N175), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[38]) );
  DFFARX1 wdata_2_reg_37_ ( .D(n808), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[37]), 
        .QN(n275) );
  DFFARX1 rdata_cp_reg_37_ ( .D(N174), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[37]) );
  DFFARX1 wdata_2_reg_36_ ( .D(n807), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[36]), 
        .QN(n274) );
  DFFARX1 rdata_cp_reg_36_ ( .D(N173), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[36]) );
  DFFARX1 wdata_2_reg_35_ ( .D(n806), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[35]), 
        .QN(n273) );
  DFFARX1 rdata_cp_reg_35_ ( .D(N172), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[35]) );
  DFFARX1 wdata_2_reg_34_ ( .D(n805), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[34]), 
        .QN(n272) );
  DFFARX1 rdata_cp_reg_34_ ( .D(N171), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[34]) );
  DFFARX1 wdata_2_reg_33_ ( .D(n804), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[33]), 
        .QN(n271) );
  DFFARX1 rdata_cp_reg_33_ ( .D(N170), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[33]) );
  DFFARX1 wdata_2_reg_32_ ( .D(n803), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[32]), 
        .QN(n270) );
  DFFARX1 rdata_cp_reg_32_ ( .D(N169), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[32]) );
  DFFARX1 wdata_2_reg_31_ ( .D(n802), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[31]), 
        .QN(n318) );
  DFFARX1 rdata_cp_reg_31_ ( .D(N168), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[31]) );
  DFFARX1 wdata_2_reg_30_ ( .D(n801), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[30]), 
        .QN(n317) );
  DFFARX1 rdata_cp_reg_30_ ( .D(N167), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[30]) );
  DFFARX1 wdata_2_reg_29_ ( .D(n800), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[29]), 
        .QN(n316) );
  DFFARX1 rdata_cp_reg_29_ ( .D(N166), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[29]) );
  DFFARX1 wdata_2_reg_28_ ( .D(n799), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[28]), 
        .QN(n315) );
  DFFARX1 rdata_cp_reg_28_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[28]) );
  DFFARX1 wdata_2_reg_27_ ( .D(n798), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[27]), 
        .QN(n314) );
  DFFARX1 rdata_cp_reg_27_ ( .D(N164), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[27]) );
  DFFARX1 wdata_2_reg_26_ ( .D(n797), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[26]), 
        .QN(n313) );
  DFFARX1 rdata_cp_reg_26_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[26]) );
  DFFARX1 wdata_2_reg_25_ ( .D(n796), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[25]), 
        .QN(n312) );
  DFFARX1 rdata_cp_reg_25_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[25]) );
  DFFARX1 wdata_2_reg_24_ ( .D(n795), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[24]), 
        .QN(n311) );
  DFFARX1 rdata_cp_reg_24_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[24]) );
  DFFARX1 wdata_2_reg_23_ ( .D(n794), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[23]), 
        .QN(n310) );
  DFFARX1 rdata_cp_reg_23_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[23]) );
  DFFARX1 wdata_2_reg_22_ ( .D(n793), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[22]), 
        .QN(n309) );
  DFFARX1 rdata_cp_reg_22_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[22]) );
  DFFARX1 wdata_2_reg_21_ ( .D(n792), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[21]), 
        .QN(n308) );
  DFFARX1 rdata_cp_reg_21_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[21]) );
  DFFARX1 wdata_2_reg_20_ ( .D(n791), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[20]), 
        .QN(n307) );
  DFFARX1 rdata_cp_reg_20_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[20]) );
  DFFARX1 wdata_2_reg_19_ ( .D(n790), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[19]), 
        .QN(n306) );
  DFFARX1 rdata_cp_reg_19_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[19]) );
  DFFARX1 wdata_2_reg_18_ ( .D(n789), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[18]), 
        .QN(n305) );
  DFFARX1 rdata_cp_reg_18_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[18]) );
  DFFARX1 wdata_2_reg_17_ ( .D(n788), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[17]), 
        .QN(n304) );
  DFFARX1 rdata_cp_reg_17_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[17]) );
  DFFARX1 wdata_2_reg_16_ ( .D(n787), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[16]), 
        .QN(n303) );
  DFFARX1 rdata_cp_reg_16_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[16]) );
  DFFARX1 wdata_2_reg_15_ ( .D(n786), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[15]), 
        .QN(n269) );
  DFFARX1 rdata_cp_reg_15_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[15]) );
  DFFARX1 wdata_2_reg_14_ ( .D(n785), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[14]), 
        .QN(n268) );
  DFFARX1 rdata_cp_reg_14_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[14]) );
  DFFARX1 wdata_2_reg_13_ ( .D(n784), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[13]), 
        .QN(n267) );
  DFFARX1 rdata_cp_reg_13_ ( .D(N150), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[13]) );
  DFFARX1 wdata_2_reg_12_ ( .D(n783), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[12]), 
        .QN(n266) );
  DFFARX1 rdata_cp_reg_12_ ( .D(N149), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[12]) );
  DFFARX1 wdata_2_reg_11_ ( .D(n782), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[11]), 
        .QN(n265) );
  DFFARX1 rdata_cp_reg_11_ ( .D(N148), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[11]) );
  DFFARX1 wdata_2_reg_10_ ( .D(n781), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[10]), 
        .QN(n264) );
  DFFARX1 rdata_cp_reg_10_ ( .D(N147), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_cp[10]) );
  DFFARX1 wdata_2_reg_9_ ( .D(n780), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[9]), 
        .QN(n302) );
  DFFARX1 rdata_cp_reg_9_ ( .D(N146), .CLK(clk), .RSTB(rst_n), .Q(rdata_cp[9])
         );
  DFFARX1 wdata_2_reg_8_ ( .D(n779), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[8]), 
        .QN(n301) );
  DFFARX1 rdata_cp_reg_8_ ( .D(N145), .CLK(clk), .RSTB(rst_n), .Q(rdata_cp[8])
         );
  DFFARX1 wdata_2_reg_7_ ( .D(n778), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[7]), 
        .QN(n326) );
  DFFARX1 wdata_2_reg_6_ ( .D(n777), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[6]), 
        .QN(n325) );
  DFFARX1 wdata_2_reg_5_ ( .D(n776), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[5]), 
        .QN(n324) );
  DFFARX1 wdata_2_reg_4_ ( .D(n775), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[4]), 
        .QN(n323) );
  DFFARX1 wdata_2_reg_3_ ( .D(n774), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[3]), 
        .QN(n322) );
  DFFARX1 wdata_2_reg_2_ ( .D(n773), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[2]), 
        .QN(n321) );
  DFFARX1 wdata_2_reg_1_ ( .D(n772), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[1]), 
        .QN(n320) );
  DFFARX1 wdata_2_reg_0_ ( .D(n771), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[0]), 
        .QN(n319) );
  DFFARX1 error_reg ( .D(n770), .CLK(clk), .RSTB(rst_n), .Q(error), .QN(n254)
         );
  XOR2X1 DP_OP_350_296_6706_U21 ( .IN1(DP_OP_350_296_6706_n40), .IN2(
        RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_1), .Q(DP_OP_350_296_6706_n22) );
  XOR2X1 DP_OP_350_296_6706_U20 ( .IN1(DP_OP_350_296_6706_n40), .IN2(
        RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_2), .Q(DP_OP_350_296_6706_n21) );
  FADDX1 DP_OP_350_296_6706_U16 ( .A(DP_OP_350_296_6706_n16), .B(address_2[1]), 
        .CI(DP_OP_350_296_6706_n22), .CO(DP_OP_350_296_6706_n15), .S(
        C36_DATA3_1) );
  FADDX1 DP_OP_350_296_6706_U15 ( .A(DP_OP_350_296_6706_n15), .B(address_2[2]), 
        .CI(DP_OP_350_296_6706_n21), .CO(DP_OP_350_296_6706_n14), .S(
        C36_DATA3_2) );
  FADDX1 DP_OP_350_296_6706_U14 ( .A(DP_OP_350_296_6706_n14), .B(address_2[3]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n13), .S(
        C36_DATA3_3) );
  FADDX1 DP_OP_350_296_6706_U13 ( .A(DP_OP_350_296_6706_n13), .B(address_2[4]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n12), .S(
        C36_DATA3_4) );
  FADDX1 DP_OP_350_296_6706_U12 ( .A(DP_OP_350_296_6706_n12), .B(address_2[5]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n11), .S(
        C36_DATA3_5) );
  FADDX1 DP_OP_350_296_6706_U11 ( .A(DP_OP_350_296_6706_n11), .B(address_2[6]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n10), .S(
        C36_DATA3_6) );
  FADDX1 DP_OP_350_296_6706_U10 ( .A(DP_OP_350_296_6706_n10), .B(address_2[7]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n9), .S(
        C36_DATA3_7) );
  FADDX1 DP_OP_350_296_6706_U9 ( .A(DP_OP_350_296_6706_n9), .B(address_2[8]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n8), .S(
        C36_DATA3_8) );
  FADDX1 DP_OP_350_296_6706_U8 ( .A(DP_OP_350_296_6706_n8), .B(address_2[9]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n7), .S(
        C36_DATA3_9) );
  FADDX1 DP_OP_350_296_6706_U7 ( .A(DP_OP_350_296_6706_n7), .B(address_2[10]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n6), .S(
        C36_DATA3_10) );
  FADDX1 DP_OP_350_296_6706_U6 ( .A(DP_OP_350_296_6706_n6), .B(address_2[11]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n5), .S(
        C36_DATA3_11) );
  FADDX1 DP_OP_350_296_6706_U5 ( .A(DP_OP_350_296_6706_n5), .B(address_2[12]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n4), .S(
        C36_DATA3_12) );
  FADDX1 DP_OP_350_296_6706_U4 ( .A(DP_OP_350_296_6706_n4), .B(address_2[13]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n3), .S(
        C36_DATA3_13) );
  FADDX1 DP_OP_350_296_6706_U3 ( .A(DP_OP_350_296_6706_n3), .B(address_2[14]), 
        .CI(DP_OP_350_296_6706_n40), .CO(DP_OP_350_296_6706_n2), .S(
        C36_DATA3_14) );
  DFFASX1 write_read_1_reg ( .D(n913), .CLK(clk), .SETB(rst_n), .Q(n203), .QN(
        n256) );
  NAND2X0 U3 ( .IN1(n914), .IN2(n913), .QN(n915) );
  NOR2X0 U4 ( .IN1(n576), .IN2(n577), .QN(n1) );
  NAND3X0 U5 ( .IN1(n579), .IN2(n578), .IN3(n1), .QN(n611) );
  XNOR2X1 U6 ( .IN1(n4), .IN2(address_2[0]), .Q(C36_DATA3_0) );
  NOR2X0 U7 ( .IN1(n559), .IN2(n560), .QN(n2) );
  NAND3X0 U8 ( .IN1(n562), .IN2(n561), .IN3(n2), .QN(n591) );
  INVX0 U9 ( .IN(counter[5]), .QN(n3) );
  NOR3X0 U10 ( .IN1(n891), .IN2(n536), .IN3(n3), .QN(n353) );
  OA21X1 U11 ( .IN1(n344), .IN2(n347), .IN3(n348), .Q(n4) );
  MUX21X1 U12 ( .IN1(address_2[0]), .IN2(DP_OP_350_296_6706_n40), .S(n4), .Q(
        DP_OP_350_296_6706_n16) );
  AOI22X1 U13 ( .IN1(n697), .IN2(n696), .IN3(n698), .IN4(n699), .QN(n5) );
  OA22X1 U14 ( .IN1(n713), .IN2(n718), .IN3(n719), .IN4(n712), .Q(n6) );
  OA22X1 U15 ( .IN1(n714), .IN2(n715), .IN3(n716), .IN4(n717), .Q(n7) );
  AND3X1 U16 ( .IN1(n5), .IN2(n6), .IN3(n7), .Q(n8) );
  NAND2X0 U17 ( .IN1(n705), .IN2(n706), .QN(n9) );
  AND2X1 U18 ( .IN1(n708), .IN2(n707), .Q(n83) );
  OA22X1 U19 ( .IN1(n883), .IN2(n675), .IN3(n736), .IN4(n887), .Q(n84) );
  NOR2X0 U20 ( .IN1(n710), .IN2(n700), .QN(n85) );
  OA22X1 U21 ( .IN1(n883), .IN2(n671), .IN3(n735), .IN4(n711), .Q(n86) );
  OA222X1 U22 ( .IN1(n9), .IN2(n83), .IN3(n84), .IN4(n85), .IN5(n86), .IN6(
        n717), .Q(n87) );
  OA22X1 U23 ( .IN1(n747), .IN2(n8), .IN3(n718), .IN4(n87), .Q(n88) );
  NOR2X0 U24 ( .IN1(n673), .IN2(n672), .QN(n89) );
  NAND3X0 U25 ( .IN1(n89), .IN2(n86), .IN3(n84), .QN(n90) );
  NOR2X0 U26 ( .IN1(n883), .IN2(n670), .QN(n91) );
  NAND4X0 U27 ( .IN1(error), .IN2(n746), .IN3(n745), .IN4(n744), .QN(n92) );
  NOR2X0 U28 ( .IN1(n91), .IN2(n92), .QN(n93) );
  NAND4X0 U29 ( .IN1(n94), .IN2(n896), .IN3(n93), .IN4(n747), .QN(n95) );
  MUX21X1 U30 ( .IN1(n301), .IN2(wdata_2[8]), .S(rdata_cp[8]), .Q(n96) );
  MUX21X1 U31 ( .IN1(n302), .IN2(wdata_2[9]), .S(rdata_cp[9]), .Q(n97) );
  MUX21X1 U32 ( .IN1(n264), .IN2(wdata_2[10]), .S(rdata_cp[10]), .Q(n98) );
  MUX21X1 U33 ( .IN1(n265), .IN2(wdata_2[11]), .S(rdata_cp[11]), .Q(n100) );
  NAND4X0 U34 ( .IN1(n96), .IN2(n97), .IN3(n98), .IN4(n100), .QN(n102) );
  MUX21X1 U35 ( .IN1(n266), .IN2(wdata_2[12]), .S(rdata_cp[12]), .Q(n104) );
  MUX21X1 U36 ( .IN1(n267), .IN2(wdata_2[13]), .S(rdata_cp[13]), .Q(n106) );
  MUX21X1 U37 ( .IN1(n268), .IN2(wdata_2[14]), .S(rdata_cp[14]), .Q(n107) );
  MUX21X1 U38 ( .IN1(n269), .IN2(wdata_2[15]), .S(rdata_cp[15]), .Q(n109) );
  NAND4X0 U39 ( .IN1(n104), .IN2(n106), .IN3(n107), .IN4(n109), .QN(n111) );
  MUX21X1 U40 ( .IN1(n303), .IN2(wdata_2[16]), .S(rdata_cp[16]), .Q(n112) );
  MUX21X1 U41 ( .IN1(n304), .IN2(wdata_2[17]), .S(rdata_cp[17]), .Q(n113) );
  MUX21X1 U42 ( .IN1(n305), .IN2(wdata_2[18]), .S(rdata_cp[18]), .Q(n116) );
  MUX21X1 U43 ( .IN1(n306), .IN2(wdata_2[19]), .S(rdata_cp[19]), .Q(n117) );
  NAND4X0 U44 ( .IN1(n112), .IN2(n113), .IN3(n116), .IN4(n117), .QN(n119) );
  MUX21X1 U45 ( .IN1(n307), .IN2(wdata_2[20]), .S(rdata_cp[20]), .Q(n120) );
  MUX21X1 U46 ( .IN1(n308), .IN2(wdata_2[21]), .S(rdata_cp[21]), .Q(n121) );
  MUX21X1 U47 ( .IN1(n309), .IN2(wdata_2[22]), .S(rdata_cp[22]), .Q(n122) );
  MUX21X1 U48 ( .IN1(n310), .IN2(wdata_2[23]), .S(rdata_cp[23]), .Q(n123) );
  NAND4X0 U49 ( .IN1(n120), .IN2(n121), .IN3(n122), .IN4(n123), .QN(n124) );
  NOR4X0 U50 ( .IN1(n102), .IN2(n111), .IN3(n119), .IN4(n124), .QN(n125) );
  MUX21X1 U51 ( .IN1(n311), .IN2(wdata_2[24]), .S(rdata_cp[24]), .Q(n126) );
  MUX21X1 U52 ( .IN1(n312), .IN2(wdata_2[25]), .S(rdata_cp[25]), .Q(n127) );
  MUX21X1 U53 ( .IN1(n313), .IN2(wdata_2[26]), .S(rdata_cp[26]), .Q(n128) );
  MUX21X1 U54 ( .IN1(n314), .IN2(wdata_2[27]), .S(rdata_cp[27]), .Q(n129) );
  NAND4X0 U55 ( .IN1(n126), .IN2(n127), .IN3(n128), .IN4(n129), .QN(n130) );
  MUX21X1 U56 ( .IN1(n315), .IN2(wdata_2[28]), .S(rdata_cp[28]), .Q(n131) );
  MUX21X1 U57 ( .IN1(n316), .IN2(wdata_2[29]), .S(rdata_cp[29]), .Q(n132) );
  MUX21X1 U58 ( .IN1(n317), .IN2(wdata_2[30]), .S(rdata_cp[30]), .Q(n133) );
  MUX21X1 U59 ( .IN1(n318), .IN2(wdata_2[31]), .S(rdata_cp[31]), .Q(n134) );
  NAND4X0 U60 ( .IN1(n131), .IN2(n132), .IN3(n133), .IN4(n134), .QN(n135) );
  MUX21X1 U61 ( .IN1(n270), .IN2(wdata_2[32]), .S(rdata_cp[32]), .Q(n136) );
  MUX21X1 U62 ( .IN1(n271), .IN2(wdata_2[33]), .S(rdata_cp[33]), .Q(n137) );
  MUX21X1 U63 ( .IN1(n272), .IN2(wdata_2[34]), .S(rdata_cp[34]), .Q(n138) );
  MUX21X1 U64 ( .IN1(n273), .IN2(wdata_2[35]), .S(rdata_cp[35]), .Q(n139) );
  NAND4X0 U65 ( .IN1(n136), .IN2(n137), .IN3(n138), .IN4(n139), .QN(n140) );
  MUX21X1 U66 ( .IN1(n274), .IN2(wdata_2[36]), .S(rdata_cp[36]), .Q(n141) );
  MUX21X1 U67 ( .IN1(n275), .IN2(wdata_2[37]), .S(rdata_cp[37]), .Q(n142) );
  MUX21X1 U68 ( .IN1(n276), .IN2(wdata_2[38]), .S(rdata_cp[38]), .Q(n143) );
  MUX21X1 U69 ( .IN1(n277), .IN2(wdata_2[39]), .S(rdata_cp[39]), .Q(n144) );
  NAND4X0 U70 ( .IN1(n141), .IN2(n142), .IN3(n143), .IN4(n144), .QN(n145) );
  NOR4X0 U71 ( .IN1(n130), .IN2(n135), .IN3(n140), .IN4(n145), .QN(n146) );
  MUX21X1 U72 ( .IN1(n278), .IN2(wdata_2[40]), .S(rdata_cp[40]), .Q(n147) );
  NAND4X0 U73 ( .IN1(n147), .IN2(n750), .IN3(n749), .IN4(n748), .QN(n148) );
  NAND4X0 U74 ( .IN1(n852), .IN2(n753), .IN3(n752), .IN4(n751), .QN(n149) );
  NAND4X0 U75 ( .IN1(n856), .IN2(n855), .IN3(n854), .IN4(n853), .QN(n150) );
  NAND4X0 U76 ( .IN1(n860), .IN2(n859), .IN3(n858), .IN4(n857), .QN(n151) );
  NOR4X0 U77 ( .IN1(n148), .IN2(n149), .IN3(n150), .IN4(n151), .QN(n152) );
  NAND4X0 U78 ( .IN1(n864), .IN2(n863), .IN3(n862), .IN4(n861), .QN(n153) );
  NAND4X0 U79 ( .IN1(n868), .IN2(n867), .IN3(n866), .IN4(n865), .QN(n154) );
  NAND4X0 U80 ( .IN1(n872), .IN2(n871), .IN3(n870), .IN4(n869), .QN(n155) );
  NAND4X0 U81 ( .IN1(n876), .IN2(n875), .IN3(n874), .IN4(n873), .QN(n156) );
  NOR4X0 U82 ( .IN1(n153), .IN2(n154), .IN3(n155), .IN4(n156), .QN(n157) );
  AND4X1 U83 ( .IN1(n125), .IN2(n146), .IN3(n152), .IN4(n157), .Q(n158) );
  NOR2X0 U84 ( .IN1(n878), .IN2(n877), .QN(n159) );
  OA22X1 U85 ( .IN1(n881), .IN2(n159), .IN3(n879), .IN4(n880), .Q(n160) );
  AOI22X1 U86 ( .IN1(n895), .IN2(n894), .IN3(n893), .IN4(n892), .QN(n161) );
  INVX0 U87 ( .IN(n888), .QN(n162) );
  OA22X1 U88 ( .IN1(n890), .IN2(n889), .IN3(n891), .IN4(n162), .Q(n163) );
  OA22X1 U89 ( .IN1(n882), .IN2(n883), .IN3(counter[0]), .IN4(n884), .Q(n164)
         );
  AO222X1 U90 ( .IN1(n887), .IN2(n886), .IN3(n887), .IN4(n164), .IN5(n886), 
        .IN6(n885), .Q(n165) );
  NAND4X0 U91 ( .IN1(n160), .IN2(n161), .IN3(n163), .IN4(n165), .QN(n166) );
  MUX21X1 U92 ( .IN1(n95), .IN2(n158), .S(n166), .Q(n167) );
  OA22X1 U93 ( .IN1(n704), .IN2(n719), .IN3(n718), .IN4(n708), .Q(n168) );
  AND4X1 U94 ( .IN1(n677), .IN2(n712), .IN3(n678), .IN4(n676), .Q(n169) );
  OA22X1 U95 ( .IN1(n714), .IN2(n169), .IN3(n716), .IN4(n85), .Q(n170) );
  AND3X1 U96 ( .IN1(n5), .IN2(n168), .IN3(n170), .Q(n171) );
  NOR2X0 U97 ( .IN1(n746), .IN2(n171), .QN(n172) );
  OAI222X1 U98 ( .IN1(n704), .IN2(n84), .IN3(n89), .IN4(n707), .IN5(n86), 
        .IN6(n712), .QN(n173) );
  INVX0 U99 ( .IN(n90), .QN(n94) );
  OA221X1 U100 ( .IN1(n173), .IN2(n697), .IN3(n173), .IN4(n90), .IN5(n701), 
        .Q(n174) );
  AOI22X1 U101 ( .IN1(n697), .IN2(n652), .IN3(n699), .IN4(n709), .QN(n175) );
  NAND3X0 U102 ( .IN1(n665), .IN2(n661), .IN3(n659), .QN(n176) );
  NAND2X0 U103 ( .IN1(n660), .IN2(n176), .QN(n177) );
  NAND2X0 U104 ( .IN1(n698), .IN2(n701), .QN(n178) );
  NAND4X0 U105 ( .IN1(n168), .IN2(n175), .IN3(n177), .IN4(n178), .QN(n179) );
  OA221X1 U106 ( .IN1(n179), .IN2(n696), .IN3(n179), .IN4(n702), .IN5(n91), 
        .Q(n180) );
  OA22X1 U107 ( .IN1(n86), .IN2(n713), .IN3(n84), .IN4(n708), .Q(n181) );
  INVX0 U108 ( .IN(n89), .QN(n182) );
  NAND3X0 U109 ( .IN1(n678), .IN2(n676), .IN3(n677), .QN(n183) );
  NAND2X0 U110 ( .IN1(n183), .IN2(n182), .QN(n184) );
  AND2X1 U111 ( .IN1(n181), .IN2(n184), .Q(n185) );
  OA22X1 U112 ( .IN1(n94), .IN2(n177), .IN3(n714), .IN4(n185), .Q(n186) );
  INVX0 U113 ( .IN(n881), .QN(n187) );
  AND3X1 U114 ( .IN1(n685), .IN2(n684), .IN3(n686), .Q(n188) );
  NAND4X0 U115 ( .IN1(n687), .IN2(n688), .IN3(n694), .IN4(n188), .QN(n189) );
  NAND4X0 U116 ( .IN1(n699), .IN2(n689), .IN3(n187), .IN4(n189), .QN(n190) );
  OR3X1 U117 ( .IN1(n84), .IN2(n719), .IN3(n169), .Q(n191) );
  AO21X1 U118 ( .IN1(n713), .IN2(n712), .IN3(n745), .Q(n192) );
  NAND4X0 U119 ( .IN1(n186), .IN2(n190), .IN3(n191), .IN4(n192), .QN(n193) );
  NOR4X0 U120 ( .IN1(n172), .IN2(n174), .IN3(n180), .IN4(n193), .QN(n194) );
  OA22X1 U121 ( .IN1(n704), .IN2(n89), .IN3(n86), .IN4(n715), .Q(n195) );
  AO21X1 U122 ( .IN1(n195), .IN2(n184), .IN3(n719), .Q(n196) );
  NAND4X0 U123 ( .IN1(n88), .IN2(n167), .IN3(n194), .IN4(n196), .QN(n770) );
  OA22X1 U124 ( .IN1(n445), .IN2(address[15]), .IN3(n446), .IN4(address[13]), 
        .Q(n197) );
  AND2X1 U125 ( .IN1(n197), .IN2(n447), .Q(n198) );
  OA222X1 U126 ( .IN1(address[11]), .IN2(n445), .IN3(n446), .IN4(address[9]), 
        .IN5(n198), .IN6(n448), .Q(n449) );
  OA22X1 U127 ( .IN1(allowable_faulty[12]), .IN2(n334), .IN3(n240), .IN4(
        allowable_faulty[11]), .Q(n199) );
  OA22X1 U128 ( .IN1(allowable_faulty[14]), .IN2(n335), .IN3(n241), .IN4(
        allowable_faulty[15]), .Q(n200) );
  NOR2X0 U129 ( .IN1(n257), .IN2(allowable_faulty[13]), .QN(n201) );
  AND3X1 U130 ( .IN1(n199), .IN2(n200), .IN3(n202), .Q(n204) );
  OA22X1 U131 ( .IN1(n332), .IN2(allowable_faulty[10]), .IN3(
        allowable_faulty[9]), .IN4(n242), .Q(n205) );
  OA22X1 U132 ( .IN1(allowable_faulty[7]), .IN2(n243), .IN3(n329), .IN4(
        allowable_faulty[8]), .Q(n206) );
  OA22X1 U133 ( .IN1(n239), .IN2(allowable_faulty[1]), .IN3(n251), .IN4(
        allowable_faulty[0]), .Q(n207) );
  AO21X1 U134 ( .IN1(allowable_faulty[1]), .IN2(n239), .IN3(n207), .Q(n208) );
  AO222X1 U135 ( .IN1(n253), .IN2(allowable_faulty[2]), .IN3(n253), .IN4(n208), 
        .IN5(allowable_faulty[2]), .IN6(n208), .Q(n209) );
  AO222X1 U136 ( .IN1(n248), .IN2(allowable_faulty[3]), .IN3(n248), .IN4(n209), 
        .IN5(allowable_faulty[3]), .IN6(n209), .Q(n210) );
  AO222X1 U137 ( .IN1(n330), .IN2(allowable_faulty[4]), .IN3(n330), .IN4(n210), 
        .IN5(allowable_faulty[4]), .IN6(n210), .Q(n211) );
  AO222X1 U138 ( .IN1(n258), .IN2(allowable_faulty[5]), .IN3(n258), .IN4(n211), 
        .IN5(allowable_faulty[5]), .IN6(n211), .Q(n212) );
  OR2X1 U139 ( .IN1(n331), .IN2(allowable_faulty[6]), .Q(n213) );
  AO222X1 U140 ( .IN1(n212), .IN2(n213), .IN3(allowable_faulty[6]), .IN4(n331), 
        .IN5(n243), .IN6(allowable_faulty[7]), .Q(n214) );
  AND4X1 U141 ( .IN1(n204), .IN2(n205), .IN3(n206), .IN4(n214), .Q(n215) );
  AO22X1 U142 ( .IN1(allowable_faulty[9]), .IN2(n242), .IN3(n329), .IN4(
        allowable_faulty[8]), .Q(n216) );
  AO222X1 U143 ( .IN1(n216), .IN2(n205), .IN3(n240), .IN4(allowable_faulty[11]), .IN5(n332), .IN6(allowable_faulty[10]), .Q(n217) );
  INVX0 U144 ( .IN(n201), .QN(n202) );
  NOR2X0 U145 ( .IN1(n201), .IN2(error_counter[12]), .QN(n218) );
  AO222X1 U146 ( .IN1(n217), .IN2(n204), .IN3(allowable_faulty[12]), .IN4(n218), .IN5(n257), .IN6(allowable_faulty[13]), .Q(n219) );
  INVX0 U147 ( .IN(error_counter[14]), .QN(n220) );
  OA21X1 U148 ( .IN1(n241), .IN2(allowable_faulty[15]), .IN3(
        allowable_faulty[14]), .Q(n221) );
  AO222X1 U149 ( .IN1(n219), .IN2(n200), .IN3(n220), .IN4(n221), .IN5(
        allowable_faulty[15]), .IN6(n241), .Q(n222) );
  NOR3X0 U150 ( .IN1(n215), .IN2(error_exceed_ignore), .IN3(n222), .QN(
        force_terminate) );
  INVX0 U151 ( .IN(n415), .QN(n223) );
  OA221X1 U152 ( .IN1(address_1[5]), .IN2(n413), .IN3(address_1[5]), .IN4(n434), .IN5(n223), .Q(N260) );
  OA22X1 U153 ( .IN1(n733), .IN2(n890), .IN3(n734), .IN4(n886), .Q(n224) );
  AOI22X1 U154 ( .IN1(n737), .IN2(n877), .IN3(n894), .IN4(n741), .QN(n225) );
  NAND2X0 U155 ( .IN1(n892), .IN2(counter[7]), .QN(n226) );
  NAND3X0 U156 ( .IN1(n226), .IN2(n880), .IN3(n724), .QN(n227) );
  NAND2X0 U157 ( .IN1(n732), .IN2(n227), .QN(n228) );
  NAND4X0 U158 ( .IN1(n742), .IN2(n224), .IN3(n225), .IN4(n228), .QN(n229) );
  NOR2X0 U159 ( .IN1(n743), .IN2(n229), .QN(n896) );
  XOR3X1 U160 ( .IN1(DP_OP_350_296_6706_n40), .IN2(DP_OP_350_296_6706_n2), 
        .IN3(address_2[15]), .Q(n230) );
  AO22X1 U161 ( .IN1(n350), .IN2(n230), .IN3(address_2[15]), .IN4(n351), .Q(
        n835) );
  INVX0 U162 ( .IN(n419), .QN(n231) );
  OA221X1 U163 ( .IN1(address_1[7]), .IN2(n417), .IN3(address_1[7]), .IN4(n434), .IN5(n231), .Q(N262) );
  NAND2X0 U164 ( .IN1(n911), .IN2(error_counter[14]), .QN(n912) );
  NAND2X0 U165 ( .IN1(n909), .IN2(error_counter[12]), .QN(n910) );
  NAND2X0 U166 ( .IN1(n907), .IN2(error_counter[10]), .QN(n908) );
  NAND2X0 U167 ( .IN1(n905), .IN2(error_counter[8]), .QN(n906) );
  NAND2X0 U168 ( .IN1(n903), .IN2(error_counter[6]), .QN(n904) );
  NAND2X0 U169 ( .IN1(n901), .IN2(error_counter[4]), .QN(n902) );
  NAND2X0 U170 ( .IN1(n437), .IN2(n436), .QN(n441) );
  NAND2X0 U171 ( .IN1(n588), .IN2(n587), .QN(n621) );
  NAND2X0 U172 ( .IN1(n616), .IN2(n597), .QN(n622) );
  NAND2X0 U173 ( .IN1(n899), .IN2(error_counter[2]), .QN(n900) );
  NAND2X0 U174 ( .IN1(n617), .IN2(n616), .QN(n626) );
  NAND2X0 U175 ( .IN1(n546), .IN2(n545), .QN(n851) );
  NAND2X0 U176 ( .IN1(n449), .IN2(n339), .QN(n340) );
  NAND2X0 U177 ( .IN1(n897), .IN2(error_counter[0]), .QN(n898) );
  NAND2X0 U178 ( .IN1(n399), .IN2(address_1[14]), .QN(n401) );
  NAND2X0 U179 ( .IN1(n599), .IN2(n598), .QN(n608) );
  NAND2X0 U180 ( .IN1(n606), .IN2(n600), .QN(n574) );
  NAND2X0 U181 ( .IN1(n448), .IN2(n397), .QN(n400) );
  NAND2X0 U182 ( .IN1(n580), .IN2(n605), .QN(n612) );
  NAND2X0 U183 ( .IN1(n504), .IN2(n507), .QN(n346) );
  NAND2X0 U184 ( .IN1(n699), .IN2(n615), .QN(n587) );
  NAND2X0 U185 ( .IN1(n718), .IN2(n615), .QN(n597) );
  NAND2X0 U186 ( .IN1(n744), .IN2(n914), .QN(n370) );
  NAND2X0 U187 ( .IN1(n556), .IN2(n555), .QN(n557) );
  NAND2X0 U188 ( .IN1(n568), .IN2(n567), .QN(n615) );
  NAND2X0 U189 ( .IN1(n565), .IN2(n564), .QN(n590) );
  NAND2X0 U190 ( .IN1(n328), .IN2(n381), .QN(n382) );
  NAND2X0 U191 ( .IN1(n681), .IN2(n680), .QN(n710) );
  NAND2X0 U192 ( .IN1(n434), .IN2(n247), .QN(n436) );
  NAND2X0 U193 ( .IN1(n467), .IN2(n466), .QN(n570) );
  NAND2X0 U194 ( .IN1(n714), .IN2(n716), .QN(n652) );
  NAND2X0 U195 ( .IN1(address_1[7]), .IN2(n417), .QN(n416) );
  NAND2X0 U196 ( .IN1(n554), .IN2(n690), .QN(n478) );
  NAND2X0 U197 ( .IN1(n694), .IN2(n693), .QN(n700) );
  NAND2X0 U198 ( .IN1(n352), .IN2(n341), .QN(n347) );
  NAND2X0 U199 ( .IN1(n487), .IN2(n554), .QN(n548) );
  NAND2X0 U200 ( .IN1(counter_1[5]), .IN2(n379), .QN(n381) );
  NAND2X0 U201 ( .IN1(n554), .IN2(n553), .QN(n555) );
  NAND2X0 U202 ( .IN1(n741), .IN2(n494), .QN(n578) );
  NAND2X0 U203 ( .IN1(n678), .IN2(n669), .QN(n702) );
  NAND2X0 U204 ( .IN1(n732), .IN2(n706), .QN(n561) );
  NAND2X0 U205 ( .IN1(n665), .IN2(n694), .QN(n698) );
  NAND2X0 U206 ( .IN1(n488), .IN2(n484), .QN(n565) );
  NAND2X0 U207 ( .IN1(n552), .IN2(n878), .QN(n502) );
  NAND2X0 U208 ( .IN1(n737), .IN2(n878), .QN(n572) );
  NAND2X0 U209 ( .IN1(n878), .IN2(n553), .QN(n501) );
  NAND2X0 U210 ( .IN1(n669), .IN2(n651), .QN(n679) );
  NAND2X0 U211 ( .IN1(n736), .IN2(n735), .QN(n877) );
  NAND2X0 U212 ( .IN1(n888), .IN2(n490), .QN(n549) );
  NAND2X0 U213 ( .IN1(n488), .IN2(n487), .QN(n571) );
  NAND2X0 U214 ( .IN1(n737), .IN2(n689), .QN(n562) );
  NAND2X0 U215 ( .IN1(n552), .IN2(n498), .QN(n485) );
  NAND2X0 U216 ( .IN1(n689), .IN2(n535), .QN(n537) );
  NAND2X0 U217 ( .IN1(n725), .IN2(n232), .QN(n670) );
  NAND2X0 U218 ( .IN1(n581), .IN2(n599), .QN(n714) );
  NAND2X0 U219 ( .IN1(n599), .IN2(n609), .QN(n719) );
  NAND2X0 U220 ( .IN1(n674), .IN2(n705), .QN(n887) );
  NAND2X0 U221 ( .IN1(n732), .IN2(n727), .QN(n733) );
  NAND2X0 U222 ( .IN1(n705), .IN2(n522), .QN(n463) );
  NAND2X0 U223 ( .IN1(n553), .IN2(n486), .QN(n491) );
  NAND2X0 U224 ( .IN1(n727), .IN2(n726), .QN(n728) );
  NAND2X0 U225 ( .IN1(counter_1[3]), .IN2(n374), .QN(n378) );
  NAND2X0 U226 ( .IN1(n481), .IN2(n528), .QN(n730) );
  NAND2X0 U227 ( .IN1(n552), .IN2(n486), .QN(n579) );
  NAND2X0 U228 ( .IN1(n674), .IN2(n895), .QN(n881) );
  NAND2X0 U229 ( .IN1(address_1[5]), .IN2(n413), .QN(n412) );
  NAND2X0 U230 ( .IN1(n726), .IN2(n232), .QN(n735) );
  NAND2X0 U231 ( .IN1(n727), .IN2(n895), .QN(n711) );
  NAND2X0 U232 ( .IN1(n727), .IN2(n705), .QN(n889) );
  NAND2X0 U233 ( .IN1(n455), .IN2(n456), .QN(n343) );
  NAND2X0 U234 ( .IN1(n528), .IN2(n530), .QN(n720) );
  NAND2X0 U235 ( .IN1(n481), .IN2(n531), .QN(n738) );
  NAND2X0 U236 ( .IN1(n718), .IN2(n610), .QN(n716) );
  NAND2X0 U237 ( .IN1(n371), .IN2(n255), .QN(n389) );
  NAND2X0 U238 ( .IN1(n497), .IN2(n538), .QN(n536) );
  NAND2X0 U239 ( .IN1(memtype[2]), .IN2(n262), .QN(n394) );
  NAND2X0 U240 ( .IN1(memtype[3]), .IN2(memtype[2]), .QN(n445) );
  NAND2X0 U241 ( .IN1(memtype[0]), .IN2(memtype[1]), .QN(n387) );
  NOR2X0 U242 ( .IN1(n916), .IN2(n480), .QN(n479) );
  AO21X1 U243 ( .IN1(n352), .IN2(n343), .IN3(n346), .Q(DP_OP_350_296_6706_n40)
         );
  NOR2X0 U244 ( .IN1(n610), .IN2(n699), .QN(n599) );
  AND4X1 U245 ( .IN1(n508), .IN2(n507), .IN3(n546), .IN4(n744), .Q(n628) );
  NAND2X0 U246 ( .IN1(address_1[1]), .IN2(n405), .QN(n406) );
  NOR2X0 U247 ( .IN1(en11), .IN2(n354), .QN(n916) );
  NAND2X0 U248 ( .IN1(n203), .IN2(n913), .QN(n480) );
  NOR2X0 U249 ( .IN1(n733), .IN2(n735), .QN(n352) );
  NAND2X0 U250 ( .IN1(n388), .IN2(n256), .QN(n438) );
  INVX0 U251 ( .IN(n916), .QN(n914) );
  INVX0 U252 ( .IN(n718), .QN(n699) );
  NOR4X0 U253 ( .IN1(en1), .IN2(en13), .IN3(en16), .IN4(en4), .QN(n718) );
  NOR2X0 U254 ( .IN1(n722), .IN2(n463), .QN(n559) );
  NOR2X0 U255 ( .IN1(n519), .IN2(n471), .QN(n689) );
  NAND2X0 U256 ( .IN1(counter[8]), .IN2(n232), .QN(n471) );
  NAND2X0 U257 ( .IN1(counter[0]), .IN2(n234), .QN(n482) );
  NOR2X0 U258 ( .IN1(memtype[0]), .IN2(memtype[1]), .QN(n386) );
  NOR2X0 U259 ( .IN1(n558), .IN2(n557), .QN(n619) );
  INVX0 U260 ( .IN(n353), .QN(n744) );
  INVX0 U261 ( .IN(n438), .QN(n434) );
  NAND2X0 U262 ( .IN1(address_1[10]), .IN2(address_1[9]), .QN(n426) );
  NOR2X0 U263 ( .IN1(n906), .IN2(n242), .QN(n907) );
  NOR2X0 U264 ( .IN1(n904), .IN2(n243), .QN(n905) );
  NOR2X0 U265 ( .IN1(n902), .IN2(n258), .QN(n903) );
  NOR2X0 U266 ( .IN1(n900), .IN2(n248), .QN(n901) );
  NOR2X0 U267 ( .IN1(n239), .IN2(n898), .QN(n899) );
  NOR2X0 U268 ( .IN1(n896), .IN2(n254), .QN(n897) );
  NOR2X0 U269 ( .IN1(n499), .IN2(n670), .QN(n566) );
  INVX0 U270 ( .IN(start), .QN(n913) );
  NOR2X0 U271 ( .IN1(DP_OP_350_296_6706_n40), .IN2(n345), .QN(n348) );
  NOR4X0 U272 ( .IN1(n353), .IN2(n346), .IN3(n352), .IN4(n345), .QN(n351) );
  NOR2X0 U273 ( .IN1(n475), .IN2(n474), .QN(n505) );
  NOR2X0 U274 ( .IN1(n570), .IN2(n473), .QN(n508) );
  NOR2X0 U275 ( .IN1(n472), .IN2(n471), .QN(n488) );
  NOR2X0 U276 ( .IN1(counter[8]), .IN2(n513), .QN(n878) );
  NAND2X0 U277 ( .IN1(counter[4]), .IN2(n233), .QN(n472) );
  NOR2X0 U278 ( .IN1(n559), .IN2(n576), .QN(n507) );
  NAND2X0 U279 ( .IN1(counter[6]), .IN2(n244), .QN(n883) );
  NAND2X0 U280 ( .IN1(n531), .IN2(n238), .QN(n477) );
  NOR2X0 U281 ( .IN1(n237), .IN2(n462), .QN(n522) );
  NAND2X0 U282 ( .IN1(counter[1]), .IN2(n235), .QN(n459) );
  NAND2X0 U283 ( .IN1(counter[6]), .IN2(counter[0]), .QN(n499) );
  INVX0 U284 ( .IN(n689), .QN(n722) );
  NAND2X0 U285 ( .IN1(counter[4]), .IN2(counter[1]), .QN(n519) );
  NAND2X0 U286 ( .IN1(counter[7]), .IN2(n705), .QN(n891) );
  INVX0 U287 ( .IN(n879), .QN(n705) );
  NAND2X0 U288 ( .IN1(n234), .IN2(n244), .QN(n879) );
  NOR2X0 U289 ( .IN1(counter[3]), .IN2(n236), .QN(n538) );
  NAND2X0 U290 ( .IN1(n245), .IN2(n357), .QN(n358) );
  NAND2X0 U291 ( .IN1(counter[5]), .IN2(n362), .QN(n364) );
  OAI21X1 U292 ( .IN1(n619), .IN2(n719), .IN3(n618), .QN(n627) );
  NOR2X0 U293 ( .IN1(n670), .IN2(n482), .QN(n560) );
  NOR2X0 U294 ( .IN1(n671), .IN2(n482), .QN(n577) );
  NOR4X0 U295 ( .IN1(n434), .IN2(n404), .IN3(n403), .IN4(n402), .QN(n433) );
  NAND2X0 U296 ( .IN1(counter_1[1]), .IN2(counter_1[0]), .QN(n373) );
  NOR2X0 U297 ( .IN1(n426), .IN2(n425), .QN(n432) );
  INVX0 U298 ( .IN(n420), .QN(n425) );
  NOR2X0 U299 ( .IN1(n250), .IN2(n416), .QN(n420) );
  NOR2X0 U300 ( .IN1(n249), .IN2(n412), .QN(n417) );
  NOR2X0 U301 ( .IN1(n499), .IN2(n671), .QN(n558) );
  INVX0 U302 ( .IN(
        RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_2), .QN(n349) );
  NOR2X0 U303 ( .IN1(n469), .IN2(n468), .QN(n556) );
  NOR2X0 U304 ( .IN1(counter[2]), .IN2(n464), .QN(n690) );
  INVX0 U305 ( .IN(n883), .QN(n895) );
  INVX0 U306 ( .IN(n489), .QN(n726) );
  NAND2X0 U307 ( .IN1(counter[2]), .IN2(counter[3]), .QN(n462) );
  NOR2X0 U308 ( .IN1(counter[7]), .IN2(n459), .QN(n531) );
  INVX0 U309 ( .IN(n884), .QN(n727) );
  INVX0 U310 ( .IN(n482), .QN(n732) );
  NOR2X0 U311 ( .IN1(n482), .IN2(n465), .QN(n552) );
  NOR2X0 U312 ( .IN1(counter[5]), .IN2(n535), .QN(n530) );
  NAND2X0 U313 ( .IN1(n236), .IN2(counter[3]), .QN(n535) );
  INVX0 U314 ( .IN(n615), .QN(n617) );
  NAND4X0 U315 ( .IN1(n575), .IN2(n584), .IN3(n587), .IN4(n574), .QN(n620) );
  NAND4X0 U316 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n583), .QN(n625) );
  AO21X1 U317 ( .IN1(n569), .IN2(n597), .IN3(n599), .Q(n584) );
  NAND3X0 U318 ( .IN1(n608), .IN2(n607), .IN3(n618), .QN(n623) );
  INVX0 U319 ( .IN(n619), .QN(n598) );
  OA222X1 U320 ( .IN1(n606), .IN2(n605), .IN3(n714), .IN4(n604), .IN5(n719), 
        .IN6(n603), .Q(n618) );
  NAND3X0 U321 ( .IN1(n573), .IN2(n572), .IN3(n571), .QN(n600) );
  INVX0 U322 ( .IN(n566), .QN(n568) );
  INVX0 U323 ( .IN(n599), .QN(n606) );
  NOR4X0 U324 ( .IN1(n577), .IN2(n560), .IN3(n743), .IN4(n506), .QN(n546) );
  AO22X1 U325 ( .IN1(address_2[0]), .IN2(n351), .IN3(n350), .IN4(C36_DATA3_0), 
        .Q(n850) );
  AO22X1 U326 ( .IN1(address_2[1]), .IN2(n351), .IN3(C36_DATA3_1), .IN4(n350), 
        .Q(n849) );
  AO22X1 U327 ( .IN1(address_2[2]), .IN2(n351), .IN3(C36_DATA3_2), .IN4(n350), 
        .Q(n848) );
  AO22X1 U328 ( .IN1(address_2[3]), .IN2(n351), .IN3(C36_DATA3_3), .IN4(n350), 
        .Q(n847) );
  AO22X1 U329 ( .IN1(address_1[1]), .IN2(n480), .IN3(address_2[1]), .IN4(n479), 
        .Q(address[1]) );
  AO22X1 U330 ( .IN1(address_1[0]), .IN2(n480), .IN3(address_2[0]), .IN4(n479), 
        .Q(address[0]) );
  AO22X1 U331 ( .IN1(address_2[4]), .IN2(n351), .IN3(C36_DATA3_4), .IN4(n350), 
        .Q(n846) );
  AO22X1 U332 ( .IN1(address_2[5]), .IN2(n351), .IN3(C36_DATA3_5), .IN4(n350), 
        .Q(n845) );
  AO22X1 U333 ( .IN1(address_2[6]), .IN2(n351), .IN3(C36_DATA3_6), .IN4(n350), 
        .Q(n844) );
  AO22X1 U334 ( .IN1(address_2[7]), .IN2(n351), .IN3(C36_DATA3_7), .IN4(n350), 
        .Q(n843) );
  AO22X1 U335 ( .IN1(address_2[8]), .IN2(n351), .IN3(C36_DATA3_8), .IN4(n350), 
        .Q(n842) );
  AO22X1 U336 ( .IN1(address_2[9]), .IN2(n351), .IN3(C36_DATA3_9), .IN4(n350), 
        .Q(n841) );
  AO22X1 U337 ( .IN1(address_2[10]), .IN2(n351), .IN3(C36_DATA3_10), .IN4(n350), .Q(n840) );
  AO22X1 U338 ( .IN1(address_2[11]), .IN2(n351), .IN3(C36_DATA3_11), .IN4(n350), .Q(n839) );
  AO22X1 U339 ( .IN1(address_2[12]), .IN2(n351), .IN3(C36_DATA3_12), .IN4(n350), .Q(n838) );
  AO22X1 U340 ( .IN1(address_2[13]), .IN2(n351), .IN3(C36_DATA3_13), .IN4(n350), .Q(n837) );
  AO22X1 U341 ( .IN1(address_2[14]), .IN2(n351), .IN3(C36_DATA3_14), .IN4(n350), .Q(n836) );
  AND2X1 U342 ( .IN1(n340), .IN2(n353), .Q(
        RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_2) );
  AO22X1 U343 ( .IN1(address_1[4]), .IN2(n480), .IN3(address_2[4]), .IN4(n479), 
        .Q(address[4]) );
  AO22X1 U344 ( .IN1(address_1[7]), .IN2(n480), .IN3(address_2[7]), .IN4(n479), 
        .Q(address[7]) );
  AO22X1 U345 ( .IN1(address_1[3]), .IN2(n480), .IN3(address_2[3]), .IN4(n479), 
        .Q(address[3]) );
  AO22X1 U346 ( .IN1(address_1[2]), .IN2(n480), .IN3(address_2[2]), .IN4(n479), 
        .Q(address[2]) );
  AO22X1 U347 ( .IN1(address_1[8]), .IN2(n480), .IN3(address_2[8]), .IN4(n479), 
        .Q(address[8]) );
  AO22X1 U348 ( .IN1(address_1[6]), .IN2(n480), .IN3(address_2[6]), .IN4(n479), 
        .Q(address[6]) );
  AO22X1 U349 ( .IN1(address_1[5]), .IN2(n480), .IN3(address_2[5]), .IN4(n479), 
        .Q(address[5]) );
  AO22X1 U350 ( .IN1(address_1[12]), .IN2(n480), .IN3(address_2[12]), .IN4(
        n479), .Q(address[12]) );
  AO22X1 U351 ( .IN1(address_1[9]), .IN2(n480), .IN3(address_2[9]), .IN4(n479), 
        .Q(address[9]) );
  AO22X1 U352 ( .IN1(address_1[11]), .IN2(n480), .IN3(address_2[11]), .IN4(
        n479), .Q(address[11]) );
  AO22X1 U353 ( .IN1(address_1[10]), .IN2(n480), .IN3(address_2[10]), .IN4(
        n479), .Q(address[10]) );
  AO22X1 U354 ( .IN1(address_1[14]), .IN2(n480), .IN3(address_2[14]), .IN4(
        n479), .Q(address[14]) );
  AO22X1 U355 ( .IN1(address_1[15]), .IN2(n480), .IN3(address_2[15]), .IN4(
        n479), .Q(address[15]) );
  AO22X1 U356 ( .IN1(address_1[13]), .IN2(n480), .IN3(address_2[13]), .IN4(
        n479), .Q(address[13]) );
  NAND3X0 U357 ( .IN1(n508), .IN2(n505), .IN3(n543), .QN(n345) );
  INVX0 U358 ( .IN(n735), .QN(n554) );
  NAND3X0 U359 ( .IN1(n488), .IN2(n530), .IN3(n895), .QN(n567) );
  NAND3X0 U360 ( .IN1(n705), .IN2(n470), .IN3(n232), .QN(n564) );
  NAND3X0 U361 ( .IN1(n878), .IN2(n895), .IN3(n690), .QN(n467) );
  INVX0 U362 ( .IN(n472), .QN(n528) );
  NAND3X0 U363 ( .IN1(n238), .IN2(n235), .IN3(n233), .QN(n489) );
  NOR3X0 U364 ( .IN1(n477), .IN2(n514), .IN3(n883), .QN(n576) );
  INVX0 U365 ( .IN(n522), .QN(n514) );
  AND3X1 U366 ( .IN1(n550), .IN2(n461), .IN3(n460), .Q(n504) );
  NOR3X0 U367 ( .IN1(counter[4]), .IN2(counter[1]), .IN3(n238), .QN(n497) );
  MUX21X1 U368 ( .IN1(n421), .IN2(n423), .S(address_1[9]), .Q(N264) );
  MUX21X1 U369 ( .IN1(n427), .IN2(n430), .S(address_1[11]), .Q(N266) );
  MUX21X1 U370 ( .IN1(n439), .IN2(n441), .S(address_1[14]), .Q(N269) );
  NOR4X0 U371 ( .IN1(en3), .IN2(en15), .IN3(en14), .IN4(en2), .QN(n581) );
  NOR2X0 U372 ( .IN1(n347), .IN2(n342), .QN(
        RSOP_343_U1_mbist_decoder_1_apnpsf_decoder_1_apnpsf_datapath_1_RSOP_343_C1_Z_1) );
  INVX0 U373 ( .IN(n344), .QN(n342) );
  NOR2X0 U374 ( .IN1(n343), .IN2(n246), .QN(n341) );
  NOR4X0 U375 ( .IN1(en10), .IN2(en12), .IN3(en2), .IN4(en4), .QN(n344) );
  OR4X1 U376 ( .IN1(en15), .IN2(en5), .IN3(en13), .IN4(en7), .Q(n246) );
  AND4X1 U377 ( .IN1(address[5]), .IN2(address[6]), .IN3(address[8]), .IN4(
        address[2]), .Q(n338) );
  AND4X1 U378 ( .IN1(n338), .IN2(n450), .IN3(address[7]), .IN4(address[4]), 
        .Q(n339) );
  NAND3X0 U379 ( .IN1(n349), .IN2(n348), .IN3(n347), .QN(n350) );
  OR4X1 U380 ( .IN1(en9), .IN2(en5), .IN3(en12), .IN4(en8), .Q(n610) );
  OR4X1 U381 ( .IN1(en7), .IN2(en10), .IN3(en6), .IN4(n714), .Q(n354) );
  NOR2X0 U382 ( .IN1(counter[0]), .IN2(n370), .QN(N111) );
  INVX0 U383 ( .IN(n370), .QN(n359) );
  OA221X1 U384 ( .IN1(counter[0]), .IN2(counter[1]), .IN3(n244), .IN4(n233), 
        .IN5(n359), .Q(N112) );
  NOR2X0 U385 ( .IN1(n244), .IN2(n233), .QN(n356) );
  NAND2X0 U386 ( .IN1(counter[0]), .IN2(counter[1]), .QN(n355) );
  OA221X1 U387 ( .IN1(counter[2]), .IN2(n356), .IN3(n236), .IN4(n355), .IN5(
        n359), .Q(N113) );
  NAND4X0 U388 ( .IN1(counter[0]), .IN2(counter[1]), .IN3(counter[2]), .IN4(
        counter[3]), .QN(n361) );
  NAND3X0 U389 ( .IN1(counter[0]), .IN2(counter[1]), .IN3(counter[2]), .QN(
        n357) );
  AND3X1 U390 ( .IN1(n361), .IN2(n359), .IN3(n358), .Q(N114) );
  INVX0 U391 ( .IN(n361), .QN(n360) );
  OA221X1 U392 ( .IN1(counter[4]), .IN2(n360), .IN3(n235), .IN4(n361), .IN5(
        n359), .Q(N115) );
  NOR2X0 U393 ( .IN1(n235), .IN2(n361), .QN(n362) );
  NOR2X0 U394 ( .IN1(n362), .IN2(counter[5]), .QN(n363) );
  INVX0 U395 ( .IN(n364), .QN(n365) );
  NOR3X0 U396 ( .IN1(n363), .IN2(n365), .IN3(n370), .QN(N116) );
  NOR2X0 U397 ( .IN1(n234), .IN2(n364), .QN(n367) );
  NOR2X0 U398 ( .IN1(n367), .IN2(n370), .QN(n366) );
  OA21X1 U399 ( .IN1(counter[6]), .IN2(n365), .IN3(n366), .Q(N117) );
  OA222X1 U400 ( .IN1(counter[7]), .IN2(n367), .IN3(counter[7]), .IN4(n914), 
        .IN5(n366), .IN6(n232), .Q(N118) );
  NAND2X0 U401 ( .IN1(counter[7]), .IN2(n367), .QN(n368) );
  MUX21X1 U402 ( .IN1(counter[8]), .IN2(n238), .S(n368), .Q(n369) );
  NOR2X0 U403 ( .IN1(n370), .IN2(n369), .QN(N119) );
  NOR4X0 U404 ( .IN1(counter_1[7]), .IN2(counter_1[4]), .IN3(counter_1[5]), 
        .IN4(counter_1[6]), .QN(n371) );
  NOR4X0 U405 ( .IN1(counter_1[1]), .IN2(counter_1[0]), .IN3(n260), .IN4(n389), 
        .QN(n388) );
  NOR2X0 U406 ( .IN1(n203), .IN2(n388), .QN(n383) );
  INVX0 U407 ( .IN(n383), .QN(n375) );
  NOR2X0 U408 ( .IN1(counter_1[0]), .IN2(n375), .QN(N133) );
  OR2X1 U409 ( .IN1(counter_1[1]), .IN2(counter_1[0]), .Q(n372) );
  AND3X1 U410 ( .IN1(n256), .IN2(n372), .IN3(n373), .Q(N134) );
  NOR2X0 U411 ( .IN1(counter_1[2]), .IN2(n373), .QN(n390) );
  OA221X1 U412 ( .IN1(n390), .IN2(counter_1[2]), .IN3(n390), .IN4(n373), .IN5(
        n383), .Q(N135) );
  NOR2X0 U413 ( .IN1(n260), .IN2(n373), .QN(n374) );
  NOR2X0 U414 ( .IN1(n374), .IN2(counter_1[3]), .QN(n376) );
  INVX0 U415 ( .IN(n378), .QN(n377) );
  NOR3X0 U416 ( .IN1(n376), .IN2(n377), .IN3(n375), .QN(N136) );
  OA221X1 U417 ( .IN1(counter_1[4]), .IN2(n377), .IN3(n327), .IN4(n378), .IN5(
        n383), .Q(N137) );
  NOR2X0 U418 ( .IN1(n327), .IN2(n378), .QN(n379) );
  OR2X1 U419 ( .IN1(counter_1[5]), .IN2(n379), .Q(n380) );
  AND3X1 U420 ( .IN1(n381), .IN2(n383), .IN3(n380), .Q(N138) );
  NOR2X0 U421 ( .IN1(n328), .IN2(n381), .QN(n385) );
  INVX0 U422 ( .IN(n385), .QN(n384) );
  AND3X1 U423 ( .IN1(n384), .IN2(n383), .IN3(n382), .Q(N139) );
  OA221X1 U424 ( .IN1(counter_1[7]), .IN2(n385), .IN3(n337), .IN4(n384), .IN5(
        n383), .Q(N140) );
  MUX21X1 U425 ( .IN1(rdata[8]), .IN2(wdata_2[8]), .S(n386), .Q(N145) );
  MUX21X1 U426 ( .IN1(rdata[9]), .IN2(wdata_2[9]), .S(n386), .Q(N146) );
  MUX21X1 U427 ( .IN1(rdata[10]), .IN2(wdata_2[10]), .S(n386), .Q(N147) );
  MUX21X1 U428 ( .IN1(rdata[11]), .IN2(wdata_2[11]), .S(n386), .Q(N148) );
  MUX21X1 U429 ( .IN1(rdata[12]), .IN2(wdata_2[12]), .S(n386), .Q(N149) );
  MUX21X1 U430 ( .IN1(rdata[13]), .IN2(wdata_2[13]), .S(n386), .Q(N150) );
  MUX21X1 U431 ( .IN1(rdata[14]), .IN2(wdata_2[14]), .S(n386), .Q(N151) );
  MUX21X1 U432 ( .IN1(rdata[15]), .IN2(wdata_2[15]), .S(n386), .Q(N152) );
  MUX21X1 U433 ( .IN1(wdata_2[16]), .IN2(rdata[16]), .S(memtype[1]), .Q(N153)
         );
  MUX21X1 U434 ( .IN1(wdata_2[17]), .IN2(rdata[17]), .S(memtype[1]), .Q(N154)
         );
  MUX21X1 U435 ( .IN1(wdata_2[18]), .IN2(rdata[18]), .S(memtype[1]), .Q(N155)
         );
  MUX21X1 U436 ( .IN1(wdata_2[19]), .IN2(rdata[19]), .S(memtype[1]), .Q(N156)
         );
  MUX21X1 U437 ( .IN1(wdata_2[20]), .IN2(rdata[20]), .S(memtype[1]), .Q(N157)
         );
  MUX21X1 U438 ( .IN1(wdata_2[21]), .IN2(rdata[21]), .S(memtype[1]), .Q(N158)
         );
  MUX21X1 U439 ( .IN1(wdata_2[22]), .IN2(rdata[22]), .S(memtype[1]), .Q(N159)
         );
  MUX21X1 U440 ( .IN1(wdata_2[23]), .IN2(rdata[23]), .S(memtype[1]), .Q(N160)
         );
  MUX21X1 U441 ( .IN1(wdata_2[24]), .IN2(rdata[24]), .S(memtype[1]), .Q(N161)
         );
  MUX21X1 U442 ( .IN1(wdata_2[25]), .IN2(rdata[25]), .S(memtype[1]), .Q(N162)
         );
  MUX21X1 U443 ( .IN1(wdata_2[26]), .IN2(rdata[26]), .S(memtype[1]), .Q(N163)
         );
  MUX21X1 U444 ( .IN1(wdata_2[27]), .IN2(rdata[27]), .S(memtype[1]), .Q(N164)
         );
  MUX21X1 U445 ( .IN1(wdata_2[28]), .IN2(rdata[28]), .S(memtype[1]), .Q(N165)
         );
  MUX21X1 U446 ( .IN1(wdata_2[29]), .IN2(rdata[29]), .S(memtype[1]), .Q(N166)
         );
  MUX21X1 U447 ( .IN1(wdata_2[30]), .IN2(rdata[30]), .S(memtype[1]), .Q(N167)
         );
  MUX21X1 U448 ( .IN1(wdata_2[31]), .IN2(rdata[31]), .S(memtype[1]), .Q(N168)
         );
  MUX21X1 U449 ( .IN1(rdata[32]), .IN2(wdata_2[32]), .S(n387), .Q(N169) );
  MUX21X1 U450 ( .IN1(rdata[33]), .IN2(wdata_2[33]), .S(n387), .Q(N170) );
  MUX21X1 U451 ( .IN1(rdata[34]), .IN2(wdata_2[34]), .S(n387), .Q(N171) );
  MUX21X1 U452 ( .IN1(rdata[35]), .IN2(wdata_2[35]), .S(n387), .Q(N172) );
  MUX21X1 U453 ( .IN1(rdata[36]), .IN2(wdata_2[36]), .S(n387), .Q(N173) );
  MUX21X1 U454 ( .IN1(rdata[37]), .IN2(wdata_2[37]), .S(n387), .Q(N174) );
  MUX21X1 U455 ( .IN1(rdata[38]), .IN2(wdata_2[38]), .S(n387), .Q(N175) );
  MUX21X1 U456 ( .IN1(rdata[39]), .IN2(wdata_2[39]), .S(n387), .Q(N176) );
  MUX21X1 U457 ( .IN1(rdata[40]), .IN2(wdata_2[40]), .S(n387), .Q(N177) );
  MUX21X1 U458 ( .IN1(rdata[41]), .IN2(wdata_2[41]), .S(n387), .Q(N178) );
  MUX21X1 U459 ( .IN1(rdata[42]), .IN2(wdata_2[42]), .S(n387), .Q(N179) );
  MUX21X1 U460 ( .IN1(rdata[43]), .IN2(wdata_2[43]), .S(n387), .Q(N180) );
  MUX21X1 U461 ( .IN1(rdata[44]), .IN2(wdata_2[44]), .S(n387), .Q(N181) );
  MUX21X1 U462 ( .IN1(rdata[45]), .IN2(wdata_2[45]), .S(n387), .Q(N182) );
  MUX21X1 U463 ( .IN1(rdata[46]), .IN2(wdata_2[46]), .S(n387), .Q(N183) );
  MUX21X1 U464 ( .IN1(rdata[47]), .IN2(wdata_2[47]), .S(n387), .Q(N184) );
  MUX21X1 U465 ( .IN1(rdata[48]), .IN2(wdata_2[48]), .S(n387), .Q(N185) );
  MUX21X1 U466 ( .IN1(rdata[49]), .IN2(wdata_2[49]), .S(n387), .Q(N186) );
  MUX21X1 U467 ( .IN1(rdata[50]), .IN2(wdata_2[50]), .S(n387), .Q(N187) );
  MUX21X1 U468 ( .IN1(rdata[51]), .IN2(wdata_2[51]), .S(n387), .Q(N188) );
  MUX21X1 U469 ( .IN1(rdata[52]), .IN2(wdata_2[52]), .S(n387), .Q(N189) );
  MUX21X1 U470 ( .IN1(rdata[53]), .IN2(wdata_2[53]), .S(n387), .Q(N190) );
  MUX21X1 U471 ( .IN1(rdata[54]), .IN2(wdata_2[54]), .S(n387), .Q(N191) );
  MUX21X1 U472 ( .IN1(rdata[55]), .IN2(wdata_2[55]), .S(n387), .Q(N192) );
  MUX21X1 U473 ( .IN1(rdata[56]), .IN2(wdata_2[56]), .S(n387), .Q(N193) );
  MUX21X1 U474 ( .IN1(rdata[57]), .IN2(wdata_2[57]), .S(n387), .Q(N194) );
  MUX21X1 U475 ( .IN1(rdata[58]), .IN2(wdata_2[58]), .S(n387), .Q(N195) );
  MUX21X1 U476 ( .IN1(rdata[59]), .IN2(wdata_2[59]), .S(n387), .Q(N196) );
  MUX21X1 U477 ( .IN1(rdata[60]), .IN2(wdata_2[60]), .S(n387), .Q(N197) );
  MUX21X1 U478 ( .IN1(rdata[61]), .IN2(wdata_2[61]), .S(n387), .Q(N198) );
  MUX21X1 U479 ( .IN1(rdata[62]), .IN2(wdata_2[62]), .S(n387), .Q(N199) );
  MUX21X1 U480 ( .IN1(rdata[63]), .IN2(wdata_2[63]), .S(n387), .Q(N200) );
  INVX0 U481 ( .IN(n389), .QN(n391) );
  NAND4X0 U482 ( .IN1(address_1[2]), .IN2(address_1[1]), .IN3(address_1[0]), 
        .IN4(address_1[3]), .QN(n409) );
  NOR2X0 U483 ( .IN1(n252), .IN2(n409), .QN(n413) );
  NAND3X0 U484 ( .IN1(n391), .IN2(n420), .IN3(n390), .QN(n392) );
  NOR2X0 U485 ( .IN1(n426), .IN2(n392), .QN(n397) );
  NAND3X0 U486 ( .IN1(address_1[11]), .IN2(address_1[12]), .IN3(n397), .QN(
        n398) );
  INVX0 U487 ( .IN(memtype[4]), .QN(n448) );
  INVX0 U488 ( .IN(n392), .QN(n393) );
  NAND3X0 U489 ( .IN1(n394), .IN2(n448), .IN3(n393), .QN(n395) );
  OA221X1 U490 ( .IN1(n398), .IN2(memtype[2]), .IN3(n398), .IN4(n247), .IN5(
        n395), .Q(n396) );
  NOR2X0 U491 ( .IN1(memtype[3]), .IN2(n396), .QN(n404) );
  NOR2X0 U492 ( .IN1(n259), .IN2(n400), .QN(n403) );
  NOR2X0 U493 ( .IN1(n247), .IN2(n398), .QN(n399) );
  OAI222X1 U494 ( .IN1(n401), .IN2(memtype[2]), .IN3(n401), .IN4(n333), .IN5(
        memtype[2]), .IN6(n400), .QN(n402) );
  MUX21X1 U495 ( .IN1(n434), .IN2(n433), .S(address_1[0]), .Q(N255) );
  NOR2X0 U496 ( .IN1(n261), .IN2(n438), .QN(n407) );
  NOR2X0 U497 ( .IN1(n433), .IN2(n261), .QN(n405) );
  OA21X1 U498 ( .IN1(address_1[1]), .IN2(n407), .IN3(n406), .Q(N256) );
  OA222X1 U499 ( .IN1(address_1[2]), .IN2(address_1[1]), .IN3(address_1[2]), 
        .IN4(n407), .IN5(n336), .IN6(n406), .Q(N257) );
  NAND3X0 U500 ( .IN1(address_1[2]), .IN2(address_1[1]), .IN3(address_1[0]), 
        .QN(n408) );
  NOR2X0 U501 ( .IN1(n438), .IN2(n408), .QN(n411) );
  OR2X1 U502 ( .IN1(n433), .IN2(n409), .Q(n410) );
  OA21X1 U503 ( .IN1(address_1[3]), .IN2(n411), .IN3(n410), .Q(N258) );
  OA222X1 U504 ( .IN1(address_1[4]), .IN2(address_1[3]), .IN3(address_1[4]), 
        .IN4(n411), .IN5(n252), .IN6(n410), .Q(N259) );
  NOR2X0 U505 ( .IN1(n433), .IN2(n412), .QN(n415) );
  NAND4X0 U506 ( .IN1(n434), .IN2(address_1[5]), .IN3(n413), .IN4(n249), .QN(
        n414) );
  OAI21X1 U507 ( .IN1(n415), .IN2(n249), .IN3(n414), .QN(N261) );
  NOR2X0 U508 ( .IN1(n433), .IN2(n416), .QN(n419) );
  NAND4X0 U509 ( .IN1(n434), .IN2(address_1[7]), .IN3(n417), .IN4(n250), .QN(
        n418) );
  OAI21X1 U510 ( .IN1(n419), .IN2(n250), .IN3(n418), .QN(N263) );
  NOR2X0 U511 ( .IN1(n438), .IN2(n425), .QN(n421) );
  OR2X1 U512 ( .IN1(n425), .IN2(n433), .Q(n423) );
  NOR2X0 U513 ( .IN1(address_1[9]), .IN2(n438), .QN(n424) );
  NOR4X0 U514 ( .IN1(address_1[10]), .IN2(n438), .IN3(n262), .IN4(n425), .QN(
        n422) );
  AO221X1 U515 ( .IN1(address_1[10]), .IN2(n424), .IN3(address_1[10]), .IN4(
        n423), .IN5(n422), .Q(N265) );
  INVX0 U516 ( .IN(n432), .QN(n428) );
  NOR2X0 U517 ( .IN1(n438), .IN2(n428), .QN(n427) );
  AO21X1 U518 ( .IN1(n428), .IN2(n434), .IN3(n433), .Q(n430) );
  NOR2X0 U519 ( .IN1(address_1[11]), .IN2(n438), .QN(n431) );
  NOR4X0 U520 ( .IN1(address_1[12]), .IN2(n259), .IN3(n438), .IN4(n428), .QN(
        n429) );
  AO221X1 U521 ( .IN1(address_1[12]), .IN2(n431), .IN3(address_1[12]), .IN4(
        n430), .IN5(n429), .Q(N267) );
  NAND3X0 U522 ( .IN1(address_1[11]), .IN2(address_1[12]), .IN3(n432), .QN(
        n435) );
  AOI21X1 U523 ( .IN1(n435), .IN2(n434), .IN3(n433), .QN(n437) );
  OAI22X1 U524 ( .IN1(n437), .IN2(n247), .IN3(n436), .IN4(n435), .QN(N268) );
  NOR3X0 U525 ( .IN1(n438), .IN2(n247), .IN3(n435), .QN(n439) );
  NOR2X0 U526 ( .IN1(address_1[14]), .IN2(n438), .QN(n442) );
  AND3X1 U527 ( .IN1(address_1[14]), .IN2(n439), .IN3(n333), .Q(n440) );
  AO221X1 U528 ( .IN1(address_1[15]), .IN2(n442), .IN3(address_1[15]), .IN4(
        n441), .IN5(n440), .Q(N270) );
  INVX0 U529 ( .IN(memtype[3]), .QN(n444) );
  OA21X1 U530 ( .IN1(address[10]), .IN2(n444), .IN3(address[3]), .Q(n450) );
  NOR2X0 U531 ( .IN1(memtype[3]), .IN2(memtype[2]), .QN(n446) );
  AND4X1 U532 ( .IN1(address[10]), .IN2(address[11]), .IN3(address[9]), .IN4(
        address[12]), .Q(n443) );
  OA21X1 U533 ( .IN1(n444), .IN2(address[14]), .IN3(n443), .Q(n447) );
  NAND3X0 U534 ( .IN1(n237), .IN2(n236), .IN3(n245), .QN(n884) );
  NOR4X0 U535 ( .IN1(address_2[4]), .IN2(address_2[8]), .IN3(address_2[5]), 
        .IN4(address_2[7]), .QN(n456) );
  NOR4X0 U536 ( .IN1(address_2[6]), .IN2(address_2[14]), .IN3(address_2[10]), 
        .IN4(address_2[15]), .QN(n454) );
  NOR4X0 U537 ( .IN1(address_2[13]), .IN2(address_2[12]), .IN3(address_2[11]), 
        .IN4(address_2[9]), .QN(n453) );
  NOR4X0 U538 ( .IN1(address_2[2]), .IN2(address_2[0]), .IN3(address_2[1]), 
        .IN4(address_2[3]), .QN(n452) );
  NOR4X0 U539 ( .IN1(en3), .IN2(en9), .IN3(en1), .IN4(en11), .QN(n451) );
  AND4X1 U540 ( .IN1(n454), .IN2(n453), .IN3(n452), .IN4(n451), .Q(n455) );
  NAND4X0 U541 ( .IN1(counter[4]), .IN2(counter[1]), .IN3(n530), .IN4(n238), 
        .QN(n729) );
  NOR2X0 U542 ( .IN1(counter[7]), .IN2(n729), .QN(n494) );
  INVX0 U543 ( .IN(n494), .QN(n675) );
  NAND3X0 U544 ( .IN1(counter[2]), .IN2(counter[3]), .IN3(n237), .QN(n465) );
  NOR2X0 U545 ( .IN1(n499), .IN2(n884), .QN(n553) );
  NOR2X0 U546 ( .IN1(n552), .IN2(n553), .QN(n734) );
  NAND4X0 U547 ( .IN1(n235), .IN2(n238), .IN3(counter[7]), .IN4(counter[1]), 
        .QN(n736) );
  INVX0 U548 ( .IN(n733), .QN(n484) );
  OR2X1 U549 ( .IN1(n237), .IN2(n535), .Q(n882) );
  NOR2X0 U550 ( .IN1(n499), .IN2(n882), .QN(n487) );
  NOR2X0 U551 ( .IN1(n484), .IN2(n487), .QN(n457) );
  OA222X1 U552 ( .IN1(n482), .IN2(n675), .IN3(n722), .IN4(n734), .IN5(n736), 
        .IN6(n457), .Q(n550) );
  NAND3X0 U553 ( .IN1(counter[2]), .IN2(counter[5]), .IN3(n245), .QN(n723) );
  NOR2X0 U554 ( .IN1(counter[8]), .IN2(n723), .QN(n481) );
  NAND4X0 U555 ( .IN1(counter[7]), .IN2(counter[4]), .IN3(counter[1]), .IN4(
        n481), .QN(n695) );
  NOR2X0 U556 ( .IN1(n232), .IN2(n482), .QN(n490) );
  NAND4X0 U557 ( .IN1(counter[8]), .IN2(n538), .IN3(n490), .IN4(n237), .QN(
        n458) );
  OA22X1 U558 ( .IN1(n482), .IN2(n695), .IN3(n459), .IN4(n458), .Q(n461) );
  NOR2X0 U559 ( .IN1(n499), .IN2(n465), .QN(n737) );
  NAND3X0 U560 ( .IN1(n737), .IN2(n531), .IN3(n238), .QN(n460) );
  NAND2X0 U561 ( .IN1(counter[7]), .IN2(n528), .QN(n513) );
  NAND2X0 U562 ( .IN1(counter[5]), .IN2(n245), .QN(n464) );
  INVX0 U563 ( .IN(n465), .QN(n674) );
  NAND4X0 U564 ( .IN1(counter[7]), .IN2(n497), .IN3(n674), .IN4(n705), .QN(
        n466) );
  INVX0 U565 ( .IN(n891), .QN(n893) );
  AND3X1 U566 ( .IN1(n726), .IN2(n530), .IN3(n893), .Q(n469) );
  NAND2X0 U567 ( .IN1(n232), .IN2(n238), .QN(n721) );
  NAND2X0 U568 ( .IN1(n538), .IN2(n237), .QN(n476) );
  NOR4X0 U569 ( .IN1(n472), .IN2(n721), .IN3(n476), .IN4(n883), .QN(n468) );
  NOR2X0 U570 ( .IN1(n237), .IN2(n536), .QN(n470) );
  NAND3X0 U571 ( .IN1(n878), .IN2(n705), .IN3(n522), .QN(n547) );
  NAND4X0 U572 ( .IN1(n556), .IN2(n564), .IN3(n547), .IN4(n567), .QN(n473) );
  INVX0 U573 ( .IN(n488), .QN(n886) );
  NOR3X0 U574 ( .IN1(n882), .IN2(n886), .IN3(n482), .QN(n475) );
  INVX0 U575 ( .IN(n548), .QN(n474) );
  AO221X1 U576 ( .IN1(n478), .IN2(n477), .IN3(n478), .IN4(n476), .IN5(n879), 
        .Q(n543) );
  OR2X1 U577 ( .IN1(n730), .IN2(counter[7]), .Q(n671) );
  NOR2X0 U578 ( .IN1(counter[5]), .IN2(n536), .QN(n725) );
  OA22X1 U579 ( .IN1(n734), .IN2(n735), .IN3(n482), .IN4(n738), .Q(n496) );
  NOR2X0 U580 ( .IN1(n235), .IN2(n233), .QN(n691) );
  NAND2X0 U581 ( .IN1(counter[7]), .IN2(n691), .QN(n483) );
  NOR2X0 U582 ( .IN1(n238), .IN2(n483), .QN(n498) );
  NAND4X0 U583 ( .IN1(n485), .IN2(n562), .IN3(n565), .IN4(n572), .QN(n493) );
  INVX0 U584 ( .IN(n736), .QN(n486) );
  NOR2X0 U585 ( .IN1(n882), .IN2(n489), .QN(n888) );
  NAND4X0 U586 ( .IN1(n491), .IN2(n579), .IN3(n571), .IN4(n549), .QN(n492) );
  NOR4X0 U587 ( .IN1(n566), .IN2(n558), .IN3(n493), .IN4(n492), .QN(n495) );
  NAND2X0 U588 ( .IN1(counter[8]), .IN2(n531), .QN(n890) );
  NOR2X0 U589 ( .IN1(n882), .IN2(n890), .QN(n706) );
  INVX0 U590 ( .IN(n499), .QN(n741) );
  NAND4X0 U591 ( .IN1(n496), .IN2(n495), .IN3(n561), .IN4(n578), .QN(n743) );
  NAND4X0 U592 ( .IN1(n741), .IN2(n497), .IN3(n522), .IN4(n232), .QN(n500) );
  INVX0 U593 ( .IN(n498), .QN(n885) );
  OA22X1 U594 ( .IN1(n499), .IN2(n695), .IN3(n885), .IN4(n733), .Q(n742) );
  NAND3X0 U595 ( .IN1(n501), .IN2(n500), .IN3(n742), .QN(n592) );
  NOR2X0 U596 ( .IN1(n352), .IN2(n592), .QN(n503) );
  NAND4X0 U597 ( .IN1(n505), .IN2(n504), .IN3(n503), .IN4(n502), .QN(n506) );
  AO221X1 U598 ( .IN1(n882), .IN2(counter[6]), .IN3(n882), .IN4(n884), .IN5(
        counter[7]), .Q(n518) );
  NAND4X0 U599 ( .IN1(counter[7]), .IN2(counter[6]), .IN3(n538), .IN4(n237), 
        .QN(n517) );
  NAND2X0 U600 ( .IN1(n522), .IN2(n234), .QN(n512) );
  NAND4X0 U601 ( .IN1(counter[4]), .IN2(n538), .IN3(n234), .IN4(n237), .QN(
        n510) );
  NAND2X0 U602 ( .IN1(n530), .IN2(n235), .QN(n509) );
  NAND4X0 U603 ( .IN1(counter[7]), .IN2(n510), .IN3(n233), .IN4(n509), .QN(
        n521) );
  INVX0 U604 ( .IN(n521), .QN(n511) );
  AO221X1 U605 ( .IN1(n232), .IN2(counter[4]), .IN3(n232), .IN4(n512), .IN5(
        n511), .Q(n515) );
  OA22X1 U606 ( .IN1(counter[1]), .IN2(n515), .IN3(n514), .IN4(n513), .Q(n516)
         );
  OA221X1 U607 ( .IN1(n519), .IN2(n518), .IN3(n519), .IN4(n517), .IN5(n516), 
        .Q(n527) );
  AO222X1 U608 ( .IN1(counter[5]), .IN2(counter[1]), .IN3(n237), .IN4(n236), 
        .IN5(counter[2]), .IN6(n233), .Q(n520) );
  NOR2X0 U609 ( .IN1(counter[3]), .IN2(n520), .QN(n529) );
  NAND3X0 U610 ( .IN1(counter[6]), .IN2(n529), .IN3(n232), .QN(n525) );
  NAND4X0 U611 ( .IN1(counter[7]), .IN2(n522), .IN3(n234), .IN4(n521), .QN(
        n524) );
  NAND3X0 U612 ( .IN1(counter[7]), .IN2(counter[1]), .IN3(n690), .QN(n523) );
  AND3X1 U613 ( .IN1(n525), .IN2(n524), .IN3(n523), .Q(n526) );
  AO221X1 U614 ( .IN1(n527), .IN2(counter[4]), .IN3(n527), .IN4(n526), .IN5(
        counter[0]), .Q(n542) );
  NOR2X0 U615 ( .IN1(n891), .IN2(n720), .QN(n534) );
  AND4X1 U616 ( .IN1(n232), .IN2(counter[4]), .IN3(n705), .IN4(n529), .Q(n533)
         );
  AND3X1 U617 ( .IN1(n531), .IN2(n530), .IN3(n244), .Q(n532) );
  NOR3X0 U618 ( .IN1(n534), .IN2(n533), .IN3(n532), .QN(n541) );
  OAI22X1 U619 ( .IN1(n538), .IN2(n537), .IN3(counter[7]), .IN4(n536), .QN(
        n539) );
  NAND3X0 U620 ( .IN1(n895), .IN2(counter[5]), .IN3(n539), .QN(n540) );
  OA221X1 U621 ( .IN1(counter[8]), .IN2(n542), .IN3(n238), .IN4(n541), .IN5(
        n540), .Q(n544) );
  NAND4X0 U622 ( .IN1(n628), .IN2(write_read_2), .IN3(n544), .IN4(n543), .QN(
        n545) );
  NAND4X0 U623 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(n551) );
  AO21X1 U624 ( .IN1(n552), .IN2(n554), .IN3(n551), .Q(n582) );
  NOR2X0 U625 ( .IN1(n582), .IN2(n598), .QN(n589) );
  NOR2X0 U626 ( .IN1(n592), .IN2(n591), .QN(n563) );
  OA22X1 U627 ( .IN1(n718), .IN2(n589), .IN3(n563), .IN4(n716), .Q(n575) );
  INVX0 U628 ( .IN(n590), .QN(n569) );
  INVX0 U629 ( .IN(n570), .QN(n573) );
  AO21X1 U630 ( .IN1(n628), .IN2(wdata_2[63]), .IN3(n620), .Q(n834) );
  NOR2X0 U631 ( .IN1(n591), .IN2(n611), .QN(n603) );
  OA22X1 U632 ( .IN1(n718), .IN2(n603), .IN3(n599), .IN4(n619), .Q(n586) );
  INVX0 U633 ( .IN(n591), .QN(n580) );
  NOR2X0 U634 ( .IN1(n590), .IN2(n615), .QN(n605) );
  NOR2X0 U635 ( .IN1(n592), .IN2(n612), .QN(n602) );
  INVX0 U636 ( .IN(n581), .QN(n609) );
  NOR2X0 U637 ( .IN1(n582), .IN2(n600), .QN(n604) );
  OA22X1 U638 ( .IN1(n602), .IN2(n719), .IN3(n604), .IN4(n716), .Q(n585) );
  NAND3X0 U639 ( .IN1(n718), .IN2(n609), .IN3(n600), .QN(n583) );
  INVX0 U640 ( .IN(n625), .QN(n588) );
  AO21X1 U641 ( .IN1(wdata_2[62]), .IN2(n628), .IN3(n621), .Q(n833) );
  NOR2X0 U642 ( .IN1(n589), .IN2(n719), .QN(n596) );
  INVX0 U643 ( .IN(n716), .QN(n701) );
  OA21X1 U644 ( .IN1(n598), .IN2(n611), .IN3(n701), .Q(n595) );
  AO22X1 U645 ( .IN1(n718), .IN2(n590), .IN3(n599), .IN4(n600), .Q(n594) );
  INVX0 U646 ( .IN(n714), .QN(n660) );
  AO22X1 U647 ( .IN1(n660), .IN2(n592), .IN3(n591), .IN4(n652), .Q(n593) );
  NOR4X0 U648 ( .IN1(n596), .IN2(n595), .IN3(n594), .IN4(n593), .QN(n616) );
  AO21X1 U649 ( .IN1(n628), .IN2(wdata_2[61]), .IN3(n622), .Q(n832) );
  INVX0 U650 ( .IN(n600), .QN(n601) );
  AO21X1 U651 ( .IN1(n602), .IN2(n601), .IN3(n718), .Q(n607) );
  AO21X1 U652 ( .IN1(n628), .IN2(wdata_2[60]), .IN3(n623), .Q(n831) );
  NOR3X0 U653 ( .IN1(n619), .IN2(n610), .IN3(n609), .QN(n614) );
  OA21X1 U654 ( .IN1(n612), .IN2(n611), .IN3(n660), .Q(n613) );
  OR3X1 U655 ( .IN1(n614), .IN2(n613), .IN3(n620), .Q(n624) );
  AO21X1 U656 ( .IN1(n628), .IN2(wdata_2[59]), .IN3(n624), .Q(n830) );
  AO21X1 U657 ( .IN1(n628), .IN2(wdata_2[58]), .IN3(n625), .Q(n829) );
  AO21X1 U658 ( .IN1(n628), .IN2(wdata_2[57]), .IN3(n626), .Q(n828) );
  AO21X1 U659 ( .IN1(n628), .IN2(wdata_2[56]), .IN3(n627), .Q(n827) );
  AO21X1 U660 ( .IN1(n628), .IN2(wdata_2[55]), .IN3(n620), .Q(n826) );
  AO21X1 U661 ( .IN1(n628), .IN2(wdata_2[54]), .IN3(n621), .Q(n825) );
  AO21X1 U662 ( .IN1(n628), .IN2(wdata_2[53]), .IN3(n622), .Q(n824) );
  AO21X1 U663 ( .IN1(n628), .IN2(wdata_2[52]), .IN3(n623), .Q(n823) );
  AO21X1 U664 ( .IN1(n628), .IN2(wdata_2[51]), .IN3(n624), .Q(n822) );
  AO21X1 U665 ( .IN1(n628), .IN2(wdata_2[50]), .IN3(n625), .Q(n821) );
  AO21X1 U666 ( .IN1(n628), .IN2(wdata_2[49]), .IN3(n626), .Q(n820) );
  AO21X1 U667 ( .IN1(n628), .IN2(wdata_2[48]), .IN3(n627), .Q(n819) );
  AO21X1 U668 ( .IN1(n628), .IN2(wdata_2[47]), .IN3(n620), .Q(n818) );
  AO21X1 U669 ( .IN1(n628), .IN2(wdata_2[46]), .IN3(n621), .Q(n817) );
  AO21X1 U670 ( .IN1(n628), .IN2(wdata_2[45]), .IN3(n622), .Q(n816) );
  AO21X1 U671 ( .IN1(n628), .IN2(wdata_2[44]), .IN3(n623), .Q(n815) );
  AO21X1 U672 ( .IN1(n628), .IN2(wdata_2[43]), .IN3(n624), .Q(n814) );
  AO21X1 U673 ( .IN1(n628), .IN2(wdata_2[42]), .IN3(n625), .Q(n813) );
  AO21X1 U674 ( .IN1(n628), .IN2(wdata_2[41]), .IN3(n626), .Q(n812) );
  AO21X1 U675 ( .IN1(n628), .IN2(wdata_2[40]), .IN3(n627), .Q(n811) );
  AO21X1 U676 ( .IN1(n628), .IN2(wdata_2[39]), .IN3(n620), .Q(n810) );
  AO21X1 U677 ( .IN1(n628), .IN2(wdata_2[38]), .IN3(n621), .Q(n809) );
  AO21X1 U678 ( .IN1(n628), .IN2(wdata_2[37]), .IN3(n622), .Q(n808) );
  AO21X1 U679 ( .IN1(n628), .IN2(wdata_2[36]), .IN3(n623), .Q(n807) );
  AO21X1 U680 ( .IN1(n628), .IN2(wdata_2[35]), .IN3(n624), .Q(n806) );
  AO21X1 U681 ( .IN1(n628), .IN2(wdata_2[34]), .IN3(n625), .Q(n805) );
  AO21X1 U682 ( .IN1(n628), .IN2(wdata_2[33]), .IN3(n626), .Q(n804) );
  AO21X1 U683 ( .IN1(n628), .IN2(wdata_2[32]), .IN3(n627), .Q(n803) );
  AO21X1 U684 ( .IN1(n628), .IN2(wdata_2[31]), .IN3(n620), .Q(n802) );
  AO21X1 U685 ( .IN1(n628), .IN2(wdata_2[30]), .IN3(n621), .Q(n801) );
  AO21X1 U686 ( .IN1(n628), .IN2(wdata_2[29]), .IN3(n622), .Q(n800) );
  AO21X1 U687 ( .IN1(n628), .IN2(wdata_2[28]), .IN3(n623), .Q(n799) );
  AO21X1 U688 ( .IN1(n628), .IN2(wdata_2[27]), .IN3(n624), .Q(n798) );
  AO21X1 U689 ( .IN1(n628), .IN2(wdata_2[26]), .IN3(n625), .Q(n797) );
  AO21X1 U690 ( .IN1(n628), .IN2(wdata_2[25]), .IN3(n626), .Q(n796) );
  AO21X1 U691 ( .IN1(n628), .IN2(wdata_2[24]), .IN3(n627), .Q(n795) );
  AO21X1 U692 ( .IN1(n628), .IN2(wdata_2[23]), .IN3(n620), .Q(n794) );
  AO21X1 U693 ( .IN1(n628), .IN2(wdata_2[22]), .IN3(n621), .Q(n793) );
  AO21X1 U694 ( .IN1(n628), .IN2(wdata_2[21]), .IN3(n622), .Q(n792) );
  AO21X1 U695 ( .IN1(n628), .IN2(wdata_2[20]), .IN3(n623), .Q(n791) );
  AO21X1 U696 ( .IN1(n628), .IN2(wdata_2[19]), .IN3(n624), .Q(n790) );
  AO21X1 U697 ( .IN1(n628), .IN2(wdata_2[18]), .IN3(n625), .Q(n789) );
  AO21X1 U698 ( .IN1(n628), .IN2(wdata_2[17]), .IN3(n626), .Q(n788) );
  AO21X1 U699 ( .IN1(n628), .IN2(wdata_2[16]), .IN3(n627), .Q(n787) );
  AO21X1 U700 ( .IN1(n628), .IN2(wdata_2[15]), .IN3(n620), .Q(n786) );
  AO21X1 U701 ( .IN1(n628), .IN2(wdata_2[14]), .IN3(n621), .Q(n785) );
  AO21X1 U702 ( .IN1(n628), .IN2(wdata_2[13]), .IN3(n622), .Q(n784) );
  AO21X1 U703 ( .IN1(n628), .IN2(wdata_2[12]), .IN3(n623), .Q(n783) );
  AO21X1 U704 ( .IN1(n628), .IN2(wdata_2[11]), .IN3(n624), .Q(n782) );
  AO21X1 U705 ( .IN1(n628), .IN2(wdata_2[10]), .IN3(n625), .Q(n781) );
  AO21X1 U706 ( .IN1(n628), .IN2(wdata_2[9]), .IN3(n626), .Q(n780) );
  AO21X1 U707 ( .IN1(n628), .IN2(wdata_2[8]), .IN3(n627), .Q(n779) );
  AO21X1 U708 ( .IN1(n628), .IN2(wdata_2[7]), .IN3(n620), .Q(n778) );
  AO21X1 U709 ( .IN1(n628), .IN2(wdata_2[6]), .IN3(n621), .Q(n777) );
  AO21X1 U710 ( .IN1(n628), .IN2(wdata_2[5]), .IN3(n622), .Q(n776) );
  AO21X1 U711 ( .IN1(n628), .IN2(wdata_2[4]), .IN3(n623), .Q(n775) );
  AO21X1 U712 ( .IN1(n628), .IN2(wdata_2[3]), .IN3(n624), .Q(n774) );
  AO21X1 U713 ( .IN1(n628), .IN2(wdata_2[2]), .IN3(n625), .Q(n773) );
  AO21X1 U714 ( .IN1(n628), .IN2(wdata_2[1]), .IN3(n626), .Q(n772) );
  AO21X1 U715 ( .IN1(n628), .IN2(wdata_2[0]), .IN3(n627), .Q(n771) );
  NAND4X0 U716 ( .IN1(rdata_cp[52]), .IN2(rdata_cp[60]), .IN3(rdata_cp[44]), 
        .IN4(rdata_cp[4]), .QN(n630) );
  NAND4X0 U717 ( .IN1(rdata_cp[28]), .IN2(rdata_cp[36]), .IN3(rdata_cp[12]), 
        .IN4(rdata_cp[20]), .QN(n629) );
  NOR2X0 U718 ( .IN1(n630), .IN2(n629), .QN(n686) );
  INVX0 U719 ( .IN(n686), .QN(n668) );
  OR4X1 U720 ( .IN1(rdata_cp[5]), .IN2(rdata_cp[61]), .IN3(rdata_cp[45]), 
        .IN4(rdata_cp[53]), .Q(n632) );
  OR4X1 U721 ( .IN1(rdata_cp[29]), .IN2(rdata_cp[37]), .IN3(rdata_cp[13]), 
        .IN4(rdata_cp[21]), .Q(n631) );
  NOR2X0 U722 ( .IN1(n632), .IN2(n631), .QN(n688) );
  NOR4X0 U723 ( .IN1(rdata_cp[57]), .IN2(rdata_cp[9]), .IN3(rdata_cp[41]), 
        .IN4(rdata_cp[49]), .QN(n634) );
  NOR4X0 U724 ( .IN1(rdata_cp[25]), .IN2(rdata_cp[33]), .IN3(rdata_cp[17]), 
        .IN4(rdata_cp[1]), .QN(n633) );
  AND3X1 U725 ( .IN1(n688), .IN2(n634), .IN3(n633), .Q(n669) );
  OR4X1 U726 ( .IN1(rdata_cp[56]), .IN2(rdata_cp[48]), .IN3(rdata_cp[8]), 
        .IN4(rdata_cp[40]), .Q(n636) );
  OR4X1 U727 ( .IN1(rdata_cp[0]), .IN2(rdata_cp[24]), .IN3(rdata_cp[32]), 
        .IN4(rdata_cp[16]), .Q(n635) );
  NOR2X0 U728 ( .IN1(n636), .IN2(n635), .QN(n651) );
  NOR2X0 U729 ( .IN1(n668), .IN2(n679), .QN(n708) );
  OR4X1 U730 ( .IN1(rdata_cp[7]), .IN2(rdata_cp[63]), .IN3(rdata_cp[55]), 
        .IN4(rdata_cp[47]), .Q(n638) );
  OR4X1 U731 ( .IN1(rdata_cp[15]), .IN2(rdata_cp[23]), .IN3(rdata_cp[39]), 
        .IN4(rdata_cp[31]), .Q(n637) );
  NOR2X0 U732 ( .IN1(n638), .IN2(n637), .QN(n659) );
  NOR4X0 U733 ( .IN1(rdata_cp[19]), .IN2(rdata_cp[35]), .IN3(rdata_cp[27]), 
        .IN4(rdata_cp[11]), .QN(n640) );
  NOR4X0 U734 ( .IN1(rdata_cp[59]), .IN2(rdata_cp[3]), .IN3(rdata_cp[51]), 
        .IN4(rdata_cp[43]), .QN(n639) );
  NAND3X0 U735 ( .IN1(n659), .IN2(n640), .IN3(n639), .QN(n682) );
  NAND4X0 U736 ( .IN1(rdata_cp[38]), .IN2(rdata_cp[14]), .IN3(rdata_cp[30]), 
        .IN4(rdata_cp[22]), .QN(n642) );
  NAND4X0 U737 ( .IN1(rdata_cp[54]), .IN2(rdata_cp[6]), .IN3(rdata_cp[62]), 
        .IN4(rdata_cp[46]), .QN(n641) );
  NOR2X0 U738 ( .IN1(n642), .IN2(n641), .QN(n687) );
  AND3X1 U739 ( .IN1(rdata_cp[18]), .IN2(rdata_cp[2]), .IN3(rdata_cp[26]), .Q(
        n644) );
  AND4X1 U740 ( .IN1(rdata_cp[58]), .IN2(rdata_cp[50]), .IN3(rdata_cp[42]), 
        .IN4(rdata_cp[34]), .Q(n643) );
  NAND4X0 U741 ( .IN1(rdata_cp[10]), .IN2(n687), .IN3(n644), .IN4(n643), .QN(
        n692) );
  NOR2X0 U742 ( .IN1(n682), .IN2(n692), .QN(n704) );
  INVX0 U743 ( .IN(n704), .QN(n709) );
  NAND4X0 U744 ( .IN1(rdata_cp[5]), .IN2(rdata_cp[61]), .IN3(rdata_cp[45]), 
        .IN4(rdata_cp[53]), .QN(n646) );
  NAND4X0 U745 ( .IN1(rdata_cp[29]), .IN2(rdata_cp[37]), .IN3(rdata_cp[13]), 
        .IN4(rdata_cp[21]), .QN(n645) );
  NOR2X0 U746 ( .IN1(n646), .IN2(n645), .QN(n676) );
  OR4X1 U747 ( .IN1(rdata_cp[52]), .IN2(rdata_cp[60]), .IN3(rdata_cp[44]), 
        .IN4(rdata_cp[4]), .Q(n648) );
  OR4X1 U748 ( .IN1(rdata_cp[28]), .IN2(rdata_cp[36]), .IN3(rdata_cp[12]), 
        .IN4(rdata_cp[20]), .Q(n647) );
  NOR2X0 U749 ( .IN1(n648), .IN2(n647), .QN(n681) );
  NAND4X0 U750 ( .IN1(rdata_cp[25]), .IN2(rdata_cp[33]), .IN3(rdata_cp[17]), 
        .IN4(rdata_cp[1]), .QN(n650) );
  NAND4X0 U751 ( .IN1(rdata_cp[57]), .IN2(rdata_cp[9]), .IN3(rdata_cp[41]), 
        .IN4(rdata_cp[49]), .QN(n649) );
  NOR2X0 U752 ( .IN1(n650), .IN2(n649), .QN(n677) );
  AND2X1 U753 ( .IN1(n677), .IN2(n651), .Q(n684) );
  NAND3X0 U754 ( .IN1(n676), .IN2(n681), .IN3(n684), .QN(n697) );
  OR4X1 U755 ( .IN1(rdata_cp[58]), .IN2(rdata_cp[50]), .IN3(rdata_cp[42]), 
        .IN4(rdata_cp[34]), .Q(n654) );
  OR4X1 U756 ( .IN1(rdata_cp[10]), .IN2(rdata_cp[18]), .IN3(rdata_cp[2]), 
        .IN4(rdata_cp[26]), .Q(n653) );
  NOR2X0 U757 ( .IN1(n654), .IN2(n653), .QN(n685) );
  NOR4X0 U758 ( .IN1(rdata_cp[54]), .IN2(rdata_cp[6]), .IN3(rdata_cp[62]), 
        .IN4(rdata_cp[46]), .QN(n656) );
  NOR4X0 U759 ( .IN1(rdata_cp[38]), .IN2(rdata_cp[14]), .IN3(rdata_cp[30]), 
        .IN4(rdata_cp[22]), .QN(n655) );
  NAND3X0 U760 ( .IN1(n685), .IN2(n656), .IN3(n655), .QN(n683) );
  INVX0 U761 ( .IN(n683), .QN(n665) );
  NAND4X0 U762 ( .IN1(rdata_cp[59]), .IN2(rdata_cp[3]), .IN3(rdata_cp[51]), 
        .IN4(rdata_cp[43]), .QN(n658) );
  NAND4X0 U763 ( .IN1(rdata_cp[19]), .IN2(rdata_cp[35]), .IN3(rdata_cp[27]), 
        .IN4(rdata_cp[11]), .QN(n657) );
  NOR2X0 U764 ( .IN1(n658), .IN2(n657), .QN(n661) );
  INVX0 U765 ( .IN(n661), .QN(n664) );
  NAND4X0 U766 ( .IN1(rdata_cp[15]), .IN2(rdata_cp[23]), .IN3(rdata_cp[39]), 
        .IN4(rdata_cp[31]), .QN(n663) );
  NAND4X0 U767 ( .IN1(rdata_cp[7]), .IN2(rdata_cp[63]), .IN3(rdata_cp[55]), 
        .IN4(rdata_cp[47]), .QN(n662) );
  NOR3X0 U768 ( .IN1(n664), .IN2(n663), .IN3(n662), .QN(n694) );
  INVX0 U769 ( .IN(n719), .QN(n696) );
  NAND4X0 U770 ( .IN1(rdata_cp[0]), .IN2(rdata_cp[24]), .IN3(rdata_cp[32]), 
        .IN4(rdata_cp[16]), .QN(n667) );
  NAND4X0 U771 ( .IN1(rdata_cp[56]), .IN2(rdata_cp[48]), .IN3(rdata_cp[8]), 
        .IN4(rdata_cp[40]), .QN(n666) );
  NOR3X0 U772 ( .IN1(n668), .IN2(n667), .IN3(n666), .QN(n678) );
  NOR2X0 U773 ( .IN1(n722), .IN2(n881), .QN(n673) );
  INVX0 U774 ( .IN(n706), .QN(n739) );
  NOR2X0 U775 ( .IN1(n739), .IN2(n879), .QN(n672) );
  INVX0 U776 ( .IN(n679), .QN(n680) );
  INVX0 U777 ( .IN(n710), .QN(n713) );
  NOR2X0 U778 ( .IN1(n683), .IN2(n682), .QN(n712) );
  NAND4X0 U779 ( .IN1(n691), .IN2(n690), .IN3(n232), .IN4(n238), .QN(n724) );
  OA22X1 U780 ( .IN1(n735), .IN2(n887), .IN3(n724), .IN4(n879), .Q(n745) );
  INVX0 U781 ( .IN(n692), .QN(n693) );
  INVX0 U782 ( .IN(n700), .QN(n707) );
  OA22X1 U783 ( .IN1(n885), .IN2(n889), .IN3(n695), .IN4(n883), .Q(n746) );
  INVX0 U784 ( .IN(n712), .QN(n703) );
  NOR2X0 U785 ( .IN1(n703), .IN2(n702), .QN(n715) );
  NOR2X0 U786 ( .IN1(n710), .IN2(n709), .QN(n717) );
  OA22X1 U787 ( .IN1(n736), .IN2(n711), .IN3(n738), .IN4(n879), .Q(n747) );
  OA22X1 U788 ( .IN1(n723), .IN2(n722), .IN3(n721), .IN4(n720), .Q(n880) );
  INVX0 U789 ( .IN(n725), .QN(n731) );
  NAND4X0 U790 ( .IN1(n731), .IN2(n730), .IN3(n729), .IN4(n728), .QN(n892) );
  NAND2X0 U791 ( .IN1(counter[7]), .IN2(n888), .QN(n740) );
  NAND3X0 U792 ( .IN1(n740), .IN2(n739), .IN3(n738), .QN(n894) );
  MUX21X1 U793 ( .IN1(n279), .IN2(wdata_2[41]), .S(rdata_cp[41]), .Q(n750) );
  MUX21X1 U794 ( .IN1(n280), .IN2(wdata_2[42]), .S(rdata_cp[42]), .Q(n749) );
  MUX21X1 U795 ( .IN1(n281), .IN2(wdata_2[43]), .S(rdata_cp[43]), .Q(n748) );
  MUX21X1 U796 ( .IN1(n282), .IN2(wdata_2[44]), .S(rdata_cp[44]), .Q(n852) );
  MUX21X1 U797 ( .IN1(n283), .IN2(wdata_2[45]), .S(rdata_cp[45]), .Q(n753) );
  MUX21X1 U798 ( .IN1(n284), .IN2(wdata_2[46]), .S(rdata_cp[46]), .Q(n752) );
  MUX21X1 U799 ( .IN1(n285), .IN2(wdata_2[47]), .S(rdata_cp[47]), .Q(n751) );
  MUX21X1 U800 ( .IN1(n286), .IN2(wdata_2[48]), .S(rdata_cp[48]), .Q(n856) );
  MUX21X1 U801 ( .IN1(n287), .IN2(wdata_2[49]), .S(rdata_cp[49]), .Q(n855) );
  MUX21X1 U802 ( .IN1(n288), .IN2(wdata_2[50]), .S(rdata_cp[50]), .Q(n854) );
  MUX21X1 U803 ( .IN1(n289), .IN2(wdata_2[51]), .S(rdata_cp[51]), .Q(n853) );
  MUX21X1 U804 ( .IN1(n290), .IN2(wdata_2[52]), .S(rdata_cp[52]), .Q(n860) );
  MUX21X1 U805 ( .IN1(n291), .IN2(wdata_2[53]), .S(rdata_cp[53]), .Q(n859) );
  MUX21X1 U806 ( .IN1(n292), .IN2(wdata_2[54]), .S(rdata_cp[54]), .Q(n858) );
  MUX21X1 U807 ( .IN1(n293), .IN2(wdata_2[55]), .S(rdata_cp[55]), .Q(n857) );
  MUX21X1 U808 ( .IN1(n294), .IN2(wdata_2[56]), .S(rdata_cp[56]), .Q(n864) );
  MUX21X1 U809 ( .IN1(n295), .IN2(wdata_2[57]), .S(rdata_cp[57]), .Q(n863) );
  MUX21X1 U810 ( .IN1(n296), .IN2(wdata_2[58]), .S(rdata_cp[58]), .Q(n862) );
  MUX21X1 U811 ( .IN1(n297), .IN2(wdata_2[59]), .S(rdata_cp[59]), .Q(n861) );
  MUX21X1 U812 ( .IN1(n298), .IN2(wdata_2[60]), .S(rdata_cp[60]), .Q(n868) );
  MUX21X1 U813 ( .IN1(n299), .IN2(wdata_2[61]), .S(rdata_cp[61]), .Q(n867) );
  MUX21X1 U814 ( .IN1(n263), .IN2(wdata_2[62]), .S(rdata_cp[62]), .Q(n866) );
  MUX21X1 U815 ( .IN1(n300), .IN2(wdata_2[63]), .S(rdata_cp[63]), .Q(n865) );
  MUX21X1 U816 ( .IN1(n326), .IN2(wdata_2[7]), .S(rdata_cp[7]), .Q(n872) );
  MUX21X1 U817 ( .IN1(n325), .IN2(wdata_2[6]), .S(rdata_cp[6]), .Q(n871) );
  MUX21X1 U818 ( .IN1(n324), .IN2(wdata_2[5]), .S(rdata_cp[5]), .Q(n870) );
  MUX21X1 U819 ( .IN1(n323), .IN2(wdata_2[4]), .S(rdata_cp[4]), .Q(n869) );
  MUX21X1 U820 ( .IN1(n322), .IN2(wdata_2[3]), .S(rdata_cp[3]), .Q(n876) );
  MUX21X1 U821 ( .IN1(n321), .IN2(wdata_2[2]), .S(rdata_cp[2]), .Q(n875) );
  MUX21X1 U822 ( .IN1(n320), .IN2(wdata_2[1]), .S(rdata_cp[1]), .Q(n874) );
  MUX21X1 U823 ( .IN1(n319), .IN2(wdata_2[0]), .S(rdata_cp[0]), .Q(n873) );
  MUX21X1 U824 ( .IN1(error_counter[0]), .IN2(n251), .S(n897), .Q(n769) );
  XNOR2X1 U825 ( .IN1(error_counter[1]), .IN2(n898), .Q(n768) );
  OA21X1 U826 ( .IN1(n899), .IN2(error_counter[2]), .IN3(n900), .Q(n767) );
  MUX21X1 U827 ( .IN1(n248), .IN2(error_counter[3]), .S(n900), .Q(n766) );
  OA21X1 U828 ( .IN1(n901), .IN2(error_counter[4]), .IN3(n902), .Q(n765) );
  MUX21X1 U829 ( .IN1(n258), .IN2(error_counter[5]), .S(n902), .Q(n764) );
  OA21X1 U830 ( .IN1(n903), .IN2(error_counter[6]), .IN3(n904), .Q(n763) );
  MUX21X1 U831 ( .IN1(n243), .IN2(error_counter[7]), .S(n904), .Q(n762) );
  OA21X1 U832 ( .IN1(n905), .IN2(error_counter[8]), .IN3(n906), .Q(n761) );
  MUX21X1 U833 ( .IN1(n242), .IN2(error_counter[9]), .S(n906), .Q(n760) );
  OA21X1 U834 ( .IN1(n907), .IN2(error_counter[10]), .IN3(n908), .Q(n759) );
  MUX21X1 U835 ( .IN1(n240), .IN2(error_counter[11]), .S(n908), .Q(n758) );
  NOR2X0 U836 ( .IN1(n908), .IN2(n240), .QN(n909) );
  OA21X1 U837 ( .IN1(n909), .IN2(error_counter[12]), .IN3(n910), .Q(n757) );
  MUX21X1 U838 ( .IN1(n257), .IN2(error_counter[13]), .S(n910), .Q(n756) );
  NOR2X0 U839 ( .IN1(n910), .IN2(n257), .QN(n911) );
  OA21X1 U840 ( .IN1(n911), .IN2(error_counter[14]), .IN3(n912), .Q(n755) );
  MUX21X1 U841 ( .IN1(n241), .IN2(error_counter[15]), .S(n912), .Q(n754) );
  NOR2X0 U842 ( .IN1(n319), .IN2(n915), .QN(wdata[0]) );
  NOR2X0 U843 ( .IN1(n264), .IN2(n915), .QN(wdata[10]) );
  NOR2X0 U844 ( .IN1(n265), .IN2(n915), .QN(wdata[11]) );
  NOR2X0 U845 ( .IN1(n266), .IN2(n915), .QN(wdata[12]) );
  NOR2X0 U846 ( .IN1(n267), .IN2(n915), .QN(wdata[13]) );
  NOR2X0 U847 ( .IN1(n268), .IN2(n915), .QN(wdata[14]) );
  NOR2X0 U848 ( .IN1(n269), .IN2(n915), .QN(wdata[15]) );
  NOR2X0 U849 ( .IN1(n303), .IN2(n915), .QN(wdata[16]) );
  NOR2X0 U850 ( .IN1(n304), .IN2(n915), .QN(wdata[17]) );
  NOR2X0 U851 ( .IN1(n305), .IN2(n915), .QN(wdata[18]) );
  NOR2X0 U852 ( .IN1(n306), .IN2(n915), .QN(wdata[19]) );
  NOR2X0 U853 ( .IN1(n320), .IN2(n915), .QN(wdata[1]) );
  NOR2X0 U854 ( .IN1(n307), .IN2(n915), .QN(wdata[20]) );
  NOR2X0 U855 ( .IN1(n308), .IN2(n915), .QN(wdata[21]) );
  NOR2X0 U856 ( .IN1(n309), .IN2(n915), .QN(wdata[22]) );
  NOR2X0 U857 ( .IN1(n310), .IN2(n915), .QN(wdata[23]) );
  NOR2X0 U858 ( .IN1(n311), .IN2(n915), .QN(wdata[24]) );
  NOR2X0 U859 ( .IN1(n312), .IN2(n915), .QN(wdata[25]) );
  NOR2X0 U860 ( .IN1(n313), .IN2(n915), .QN(wdata[26]) );
  NOR2X0 U861 ( .IN1(n314), .IN2(n915), .QN(wdata[27]) );
  NOR2X0 U862 ( .IN1(n315), .IN2(n915), .QN(wdata[28]) );
  NOR2X0 U863 ( .IN1(n316), .IN2(n915), .QN(wdata[29]) );
  NOR2X0 U864 ( .IN1(n321), .IN2(n915), .QN(wdata[2]) );
  NOR2X0 U865 ( .IN1(n317), .IN2(n915), .QN(wdata[30]) );
  NOR2X0 U866 ( .IN1(n318), .IN2(n915), .QN(wdata[31]) );
  NOR2X0 U867 ( .IN1(n270), .IN2(n915), .QN(wdata[32]) );
  NOR2X0 U868 ( .IN1(n271), .IN2(n915), .QN(wdata[33]) );
  NOR2X0 U869 ( .IN1(n272), .IN2(n915), .QN(wdata[34]) );
  NOR2X0 U870 ( .IN1(n273), .IN2(n915), .QN(wdata[35]) );
  NOR2X0 U871 ( .IN1(n274), .IN2(n915), .QN(wdata[36]) );
  NOR2X0 U872 ( .IN1(n275), .IN2(n915), .QN(wdata[37]) );
  NOR2X0 U873 ( .IN1(n276), .IN2(n915), .QN(wdata[38]) );
  NOR2X0 U874 ( .IN1(n277), .IN2(n915), .QN(wdata[39]) );
  NOR2X0 U875 ( .IN1(n322), .IN2(n915), .QN(wdata[3]) );
  NOR2X0 U876 ( .IN1(n278), .IN2(n915), .QN(wdata[40]) );
  NOR2X0 U877 ( .IN1(n279), .IN2(n915), .QN(wdata[41]) );
  NOR2X0 U878 ( .IN1(n280), .IN2(n915), .QN(wdata[42]) );
  NOR2X0 U879 ( .IN1(n281), .IN2(n915), .QN(wdata[43]) );
  NOR2X0 U880 ( .IN1(n282), .IN2(n915), .QN(wdata[44]) );
  NOR2X0 U881 ( .IN1(n283), .IN2(n915), .QN(wdata[45]) );
  NOR2X0 U882 ( .IN1(n284), .IN2(n915), .QN(wdata[46]) );
  NOR2X0 U883 ( .IN1(n285), .IN2(n915), .QN(wdata[47]) );
  NOR2X0 U884 ( .IN1(n286), .IN2(n915), .QN(wdata[48]) );
  NOR2X0 U885 ( .IN1(n287), .IN2(n915), .QN(wdata[49]) );
  NOR2X0 U886 ( .IN1(n323), .IN2(n915), .QN(wdata[4]) );
  NOR2X0 U887 ( .IN1(n288), .IN2(n915), .QN(wdata[50]) );
  NOR2X0 U888 ( .IN1(n289), .IN2(n915), .QN(wdata[51]) );
  NOR2X0 U889 ( .IN1(n290), .IN2(n915), .QN(wdata[52]) );
  NOR2X0 U890 ( .IN1(n291), .IN2(n915), .QN(wdata[53]) );
  NOR2X0 U891 ( .IN1(n292), .IN2(n915), .QN(wdata[54]) );
  NOR2X0 U892 ( .IN1(n293), .IN2(n915), .QN(wdata[55]) );
  NOR2X0 U893 ( .IN1(n294), .IN2(n915), .QN(wdata[56]) );
  NOR2X0 U894 ( .IN1(n295), .IN2(n915), .QN(wdata[57]) );
  NOR2X0 U895 ( .IN1(n296), .IN2(n915), .QN(wdata[58]) );
  NOR2X0 U896 ( .IN1(n297), .IN2(n915), .QN(wdata[59]) );
  NOR2X0 U897 ( .IN1(n324), .IN2(n915), .QN(wdata[5]) );
  NOR2X0 U898 ( .IN1(n298), .IN2(n915), .QN(wdata[60]) );
  NOR2X0 U899 ( .IN1(n299), .IN2(n915), .QN(wdata[61]) );
  NOR2X0 U900 ( .IN1(n263), .IN2(n915), .QN(wdata[62]) );
  NOR2X0 U901 ( .IN1(n300), .IN2(n915), .QN(wdata[63]) );
  NOR2X0 U902 ( .IN1(n325), .IN2(n915), .QN(wdata[6]) );
  NOR2X0 U903 ( .IN1(n326), .IN2(n915), .QN(wdata[7]) );
  NOR2X0 U904 ( .IN1(n301), .IN2(n915), .QN(wdata[8]) );
  NOR2X0 U905 ( .IN1(n302), .IN2(n915), .QN(wdata[9]) );
  NOR2X0 U906 ( .IN1(n916), .IN2(start), .QN(n917) );
  AO21X1 U907 ( .IN1(write_read_2), .IN2(n917), .IN3(n256), .Q(write_read) );
endmodule


module apnpsf_decoder ( clk, rst_n, apnpsf_en, error_exceed_ignore, 
        allowable_faulty, address, write_read, memtype, wdata, rdata, error, 
        force_terminate, apnpsf_complete );
  input [15:0] allowable_faulty;
  output [15:0] address;
  input [4:0] memtype;
  output [63:0] wdata;
  input [63:0] rdata;
  input clk, rst_n, apnpsf_en, error_exceed_ignore;
  output write_read, error, force_terminate, apnpsf_complete;
  wire   start, en1, en2, en3, en4, en5, en6, en7, en8, en9, en10, en11, en12,
         en13, en14, en15, en16;
  wire   [8:0] counter;

  apnpsf_controller apnpsf_controller_1 ( .clk(clk), .rst_n(rst_n), 
        .apnpsf_en(apnpsf_en), .memtype({memtype[4:2], 1'b0, 1'b0}), .address(
        address), .counter(counter), .start(start), .en1(en1), .en2(en2), 
        .en3(en3), .en4(en4), .en5(en5), .en6(en6), .en7(en7), .en8(en8), 
        .en9(en9), .en10(en10), .en11(en11), .en12(en12), .en13(en13), .en14(
        en14), .en15(en15), .en16(en16), .finish(apnpsf_complete) );
  apnpsf_datapath apnpsf_datapath_1 ( .clk(clk), .rst_n(rst_n), .start(start), 
        .en1(en1), .en2(en2), .en3(en3), .en4(en4), .en5(en5), .en6(en6), 
        .en7(en7), .en8(en8), .en9(en9), .en10(en10), .en11(en11), .en12(en12), 
        .en13(en13), .en14(en14), .en15(en15), .en16(en16), 
        .error_exceed_ignore(error_exceed_ignore), .allowable_faulty(
        allowable_faulty), .address(address), .write_read(write_read), .wdata(
        wdata), .rdata(rdata), .counter(counter), .error(error), 
        .force_terminate(force_terminate), .memtype(memtype) );
endmodule


module mbist_decoder ( clk, rst_n, apnpsf_en, error_exceed_ignore, 
        allowable_faulty, memtype, address, write_read, wdata, rdata, error, 
        force_terminate, apnpsf_complete );
  input [15:0] allowable_faulty;
  input [4:0] memtype;
  output [15:0] address;
  output [63:0] wdata;
  input [63:0] rdata;
  input clk, rst_n, apnpsf_en, error_exceed_ignore;
  output write_read, error, force_terminate, apnpsf_complete;
  wire   apnpsf_write_read, apnpsf_error, apnpsf_force_terminate, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84;
  wire   [15:0] apnpsf_address;
  wire   [63:0] apnpsf_wdata;

  apnpsf_decoder apnpsf_decoder_1 ( .clk(clk), .rst_n(rst_n), .apnpsf_en(
        apnpsf_en), .error_exceed_ignore(error_exceed_ignore), 
        .allowable_faulty(allowable_faulty), .address(apnpsf_address), 
        .write_read(apnpsf_write_read), .memtype(memtype), .wdata(apnpsf_wdata), .rdata(rdata), .error(apnpsf_error), .force_terminate(apnpsf_force_terminate), .apnpsf_complete(apnpsf_complete) );
  DFFARX1 wdata_reg_63_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(wdata[63]) );
  DFFARX1 wdata_reg_62_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(wdata[62]) );
  DFFARX1 wdata_reg_61_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(wdata[61]) );
  DFFARX1 wdata_reg_60_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(wdata[60]) );
  DFFARX1 wdata_reg_59_ ( .D(N80), .CLK(clk), .RSTB(rst_n), .Q(wdata[59]) );
  DFFARX1 wdata_reg_58_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(wdata[58]) );
  DFFARX1 wdata_reg_57_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(wdata[57]) );
  DFFARX1 wdata_reg_56_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(wdata[56]) );
  DFFARX1 wdata_reg_55_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(wdata[55]) );
  DFFARX1 wdata_reg_54_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(wdata[54]) );
  DFFARX1 wdata_reg_53_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(wdata[53]) );
  DFFARX1 wdata_reg_52_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(wdata[52]) );
  DFFARX1 wdata_reg_51_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(wdata[51]) );
  DFFARX1 wdata_reg_50_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(wdata[50]) );
  DFFARX1 wdata_reg_49_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(wdata[49]) );
  DFFARX1 wdata_reg_48_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(wdata[48]) );
  DFFARX1 wdata_reg_47_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(wdata[47]) );
  DFFARX1 wdata_reg_46_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(wdata[46]) );
  DFFARX1 wdata_reg_45_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(wdata[45]) );
  DFFARX1 wdata_reg_44_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(wdata[44]) );
  DFFARX1 wdata_reg_43_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(wdata[43]) );
  DFFARX1 wdata_reg_42_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(wdata[42]) );
  DFFARX1 wdata_reg_41_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(wdata[41]) );
  DFFARX1 wdata_reg_40_ ( .D(N61), .CLK(clk), .RSTB(rst_n), .Q(wdata[40]) );
  DFFARX1 wdata_reg_39_ ( .D(N60), .CLK(clk), .RSTB(rst_n), .Q(wdata[39]) );
  DFFARX1 wdata_reg_38_ ( .D(N59), .CLK(clk), .RSTB(rst_n), .Q(wdata[38]) );
  DFFARX1 wdata_reg_37_ ( .D(N58), .CLK(clk), .RSTB(rst_n), .Q(wdata[37]) );
  DFFARX1 wdata_reg_36_ ( .D(N57), .CLK(clk), .RSTB(rst_n), .Q(wdata[36]) );
  DFFARX1 wdata_reg_35_ ( .D(N56), .CLK(clk), .RSTB(rst_n), .Q(wdata[35]) );
  DFFARX1 wdata_reg_34_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(wdata[34]) );
  DFFARX1 wdata_reg_33_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(wdata[33]) );
  DFFARX1 wdata_reg_32_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(wdata[32]) );
  DFFARX1 wdata_reg_31_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(wdata[31]) );
  DFFARX1 wdata_reg_30_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(wdata[30]) );
  DFFARX1 wdata_reg_29_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(wdata[29]) );
  DFFARX1 wdata_reg_28_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(wdata[28]) );
  DFFARX1 wdata_reg_27_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(wdata[27]) );
  DFFARX1 wdata_reg_26_ ( .D(N47), .CLK(clk), .RSTB(rst_n), .Q(wdata[26]) );
  DFFARX1 wdata_reg_25_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(wdata[25]) );
  DFFARX1 wdata_reg_24_ ( .D(N45), .CLK(clk), .RSTB(rst_n), .Q(wdata[24]) );
  DFFARX1 wdata_reg_23_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(wdata[23]) );
  DFFARX1 wdata_reg_22_ ( .D(N43), .CLK(clk), .RSTB(rst_n), .Q(wdata[22]) );
  DFFARX1 wdata_reg_21_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(wdata[21]) );
  DFFARX1 wdata_reg_20_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(wdata[20]) );
  DFFARX1 wdata_reg_19_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(wdata[19]) );
  DFFARX1 wdata_reg_18_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(wdata[18]) );
  DFFARX1 wdata_reg_17_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(wdata[17]) );
  DFFARX1 wdata_reg_16_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(wdata[16]) );
  DFFARX1 wdata_reg_15_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(wdata[15]) );
  DFFARX1 wdata_reg_14_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(wdata[14]) );
  DFFARX1 wdata_reg_13_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(wdata[13]) );
  DFFARX1 wdata_reg_12_ ( .D(N33), .CLK(clk), .RSTB(rst_n), .Q(wdata[12]) );
  DFFARX1 wdata_reg_11_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(wdata[11]) );
  DFFARX1 wdata_reg_10_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(wdata[10]) );
  DFFARX1 wdata_reg_9_ ( .D(N30), .CLK(clk), .RSTB(rst_n), .Q(wdata[9]) );
  DFFARX1 wdata_reg_8_ ( .D(N29), .CLK(clk), .RSTB(rst_n), .Q(wdata[8]) );
  DFFARX1 wdata_reg_7_ ( .D(N28), .CLK(clk), .RSTB(rst_n), .Q(wdata[7]) );
  DFFARX1 wdata_reg_6_ ( .D(N27), .CLK(clk), .RSTB(rst_n), .Q(wdata[6]) );
  DFFARX1 wdata_reg_5_ ( .D(N26), .CLK(clk), .RSTB(rst_n), .Q(wdata[5]) );
  DFFARX1 wdata_reg_4_ ( .D(N25), .CLK(clk), .RSTB(rst_n), .Q(wdata[4]) );
  DFFARX1 wdata_reg_3_ ( .D(N24), .CLK(clk), .RSTB(rst_n), .Q(wdata[3]) );
  DFFARX1 wdata_reg_2_ ( .D(N23), .CLK(clk), .RSTB(rst_n), .Q(wdata[2]) );
  DFFARX1 wdata_reg_1_ ( .D(N22), .CLK(clk), .RSTB(rst_n), .Q(wdata[1]) );
  DFFARX1 wdata_reg_0_ ( .D(N21), .CLK(clk), .RSTB(rst_n), .Q(wdata[0]) );
  AND2X1 U3 ( .IN1(apnpsf_en), .IN2(apnpsf_write_read), .Q(write_read) );
  AND2X1 U5 ( .IN1(apnpsf_en), .IN2(apnpsf_error), .Q(error) );
  AND2X1 U22 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[63]), .Q(N84) );
  AND2X1 U23 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[62]), .Q(N83) );
  AND2X1 U24 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[61]), .Q(N82) );
  AND2X1 U25 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[60]), .Q(N81) );
  AND2X1 U26 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[59]), .Q(N80) );
  AND2X1 U27 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[58]), .Q(N79) );
  AND2X1 U28 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[57]), .Q(N78) );
  AND2X1 U29 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[56]), .Q(N77) );
  AND2X1 U30 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[55]), .Q(N76) );
  AND2X1 U31 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[54]), .Q(N75) );
  AND2X1 U32 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[53]), .Q(N74) );
  AND2X1 U33 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[52]), .Q(N73) );
  AND2X1 U34 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[51]), .Q(N72) );
  AND2X1 U35 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[50]), .Q(N71) );
  AND2X1 U36 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[49]), .Q(N70) );
  AND2X1 U37 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[48]), .Q(N69) );
  AND2X1 U38 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[47]), .Q(N68) );
  AND2X1 U39 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[46]), .Q(N67) );
  AND2X1 U40 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[45]), .Q(N66) );
  AND2X1 U41 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[44]), .Q(N65) );
  AND2X1 U42 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[43]), .Q(N64) );
  AND2X1 U43 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[42]), .Q(N63) );
  AND2X1 U44 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[41]), .Q(N62) );
  AND2X1 U45 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[40]), .Q(N61) );
  AND2X1 U46 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[39]), .Q(N60) );
  AND2X1 U47 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[38]), .Q(N59) );
  AND2X1 U48 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[37]), .Q(N58) );
  AND2X1 U49 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[36]), .Q(N57) );
  AND2X1 U50 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[35]), .Q(N56) );
  AND2X1 U51 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[34]), .Q(N55) );
  AND2X1 U52 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[33]), .Q(N54) );
  AND2X1 U53 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[32]), .Q(N53) );
  AND2X1 U54 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[31]), .Q(N52) );
  AND2X1 U55 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[30]), .Q(N51) );
  AND2X1 U56 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[29]), .Q(N50) );
  AND2X1 U57 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[28]), .Q(N49) );
  AND2X1 U58 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[27]), .Q(N48) );
  AND2X1 U59 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[26]), .Q(N47) );
  AND2X1 U60 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[25]), .Q(N46) );
  AND2X1 U61 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[24]), .Q(N45) );
  AND2X1 U62 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[23]), .Q(N44) );
  AND2X1 U63 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[22]), .Q(N43) );
  AND2X1 U64 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[21]), .Q(N42) );
  AND2X1 U65 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[20]), .Q(N41) );
  AND2X1 U66 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[19]), .Q(N40) );
  AND2X1 U67 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[18]), .Q(N39) );
  AND2X1 U68 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[17]), .Q(N38) );
  AND2X1 U69 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[16]), .Q(N37) );
  AND2X1 U70 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[15]), .Q(N36) );
  AND2X1 U71 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[14]), .Q(N35) );
  AND2X1 U72 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[13]), .Q(N34) );
  AND2X1 U73 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[12]), .Q(N33) );
  AND2X1 U74 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[11]), .Q(N32) );
  AND2X1 U75 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[10]), .Q(N31) );
  AND2X1 U76 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[9]), .Q(N30) );
  AND2X1 U77 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[8]), .Q(N29) );
  AND2X1 U78 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[7]), .Q(N28) );
  AND2X1 U79 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[6]), .Q(N27) );
  AND2X1 U80 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[5]), .Q(N26) );
  AND2X1 U81 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[4]), .Q(N25) );
  AND2X1 U82 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[3]), .Q(N24) );
  AND2X1 U83 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[2]), .Q(N23) );
  AND2X1 U84 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[1]), .Q(N22) );
  AND2X1 U85 ( .IN1(apnpsf_en), .IN2(apnpsf_wdata[0]), .Q(N21) );
  AND2X1 U11 ( .IN1(apnpsf_en), .IN2(apnpsf_address[4]), .Q(address[4]) );
  AND2X1 U10 ( .IN1(apnpsf_en), .IN2(apnpsf_address[5]), .Q(address[5]) );
  AND2X1 U9 ( .IN1(apnpsf_en), .IN2(apnpsf_address[6]), .Q(address[6]) );
  AND2X1 U8 ( .IN1(apnpsf_en), .IN2(apnpsf_address[7]), .Q(address[7]) );
  AND2X1 U7 ( .IN1(apnpsf_en), .IN2(apnpsf_address[8]), .Q(address[8]) );
  AND2X1 U6 ( .IN1(apnpsf_en), .IN2(apnpsf_address[9]), .Q(address[9]) );
  AND2X1 U20 ( .IN1(apnpsf_en), .IN2(apnpsf_address[10]), .Q(address[10]) );
  AND2X1 U19 ( .IN1(apnpsf_en), .IN2(apnpsf_address[11]), .Q(address[11]) );
  AND2X1 U18 ( .IN1(apnpsf_en), .IN2(apnpsf_address[12]), .Q(address[12]) );
  AND2X1 U17 ( .IN1(apnpsf_en), .IN2(apnpsf_address[13]), .Q(address[13]) );
  AND2X1 U16 ( .IN1(apnpsf_en), .IN2(apnpsf_address[14]), .Q(address[14]) );
  AND2X1 U15 ( .IN1(apnpsf_en), .IN2(apnpsf_address[15]), .Q(address[15]) );
  AND2X1 U14 ( .IN1(apnpsf_en), .IN2(apnpsf_address[1]), .Q(address[1]) );
  AND2X1 U13 ( .IN1(apnpsf_en), .IN2(apnpsf_address[2]), .Q(address[2]) );
  AND2X1 U12 ( .IN1(apnpsf_en), .IN2(apnpsf_address[3]), .Q(address[3]) );
  AND2X1 U21 ( .IN1(apnpsf_en), .IN2(apnpsf_address[0]), .Q(address[0]) );
  AND2X1 U4 ( .IN1(apnpsf_en), .IN2(apnpsf_force_terminate), .Q(
        force_terminate) );
endmodule


module mbist_mux_demux ( clk, rst_n, memory_sel, write_read_mbist, rdata_mbist, 
        wdata_mbist, address_mbist, write_read_7, write_read_6, write_read_5, 
        write_read_4, write_read_3, write_read_2, write_read_1, write_read_0, 
        rdata_7, rdata_6, rdata_5, rdata_4, rdata_3, rdata_2, rdata_1, rdata_0, 
        wdata_7, wdata_6, wdata_5, wdata_4, wdata_3, wdata_2, wdata_1, wdata_0, 
        address_7, address_6, address_5, address_4, address_3, address_2, 
        address_1, address_0 );
  input [2:0] memory_sel;
  output [63:0] rdata_mbist;
  input [63:0] wdata_mbist;
  input [15:0] address_mbist;
  input [63:0] rdata_7;
  input [63:0] rdata_6;
  input [63:0] rdata_5;
  input [63:0] rdata_4;
  input [63:0] rdata_3;
  input [63:0] rdata_2;
  input [63:0] rdata_1;
  input [63:0] rdata_0;
  output [63:0] wdata_7;
  output [63:0] wdata_6;
  output [63:0] wdata_5;
  output [63:0] wdata_4;
  output [63:0] wdata_3;
  output [63:0] wdata_2;
  output [63:0] wdata_1;
  output [63:0] wdata_0;
  output [15:0] address_7;
  output [15:0] address_6;
  output [15:0] address_5;
  output [15:0] address_4;
  output [15:0] address_3;
  output [15:0] address_2;
  output [15:0] address_1;
  output [15:0] address_0;
  input clk, rst_n, write_read_mbist;
  output write_read_7, write_read_6, write_read_5, write_read_4, write_read_3,
         write_read_2, write_read_1, write_read_0;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694,
         N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705,
         N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716,
         N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n713, n714, n715,
         n716, n717, n718, n719, n720;

  DFFARX1 address_4_reg_15_ ( .D(N144), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[15]) );
  DFFARX1 address_4_reg_14_ ( .D(N143), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[14]) );
  DFFARX1 address_4_reg_13_ ( .D(N142), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[13]) );
  DFFARX1 address_4_reg_12_ ( .D(N141), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[12]) );
  DFFARX1 address_4_reg_11_ ( .D(N140), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[11]) );
  DFFARX1 address_4_reg_10_ ( .D(N139), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[10]) );
  DFFARX1 address_4_reg_9_ ( .D(N138), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[9]) );
  DFFARX1 address_4_reg_8_ ( .D(N137), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[8]) );
  DFFARX1 address_4_reg_7_ ( .D(N136), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[7]) );
  DFFARX1 address_4_reg_6_ ( .D(N135), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[6]) );
  DFFARX1 address_4_reg_5_ ( .D(N134), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[5]) );
  DFFARX1 address_4_reg_4_ ( .D(N133), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[4]) );
  DFFARX1 address_4_reg_3_ ( .D(N132), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[3]) );
  DFFARX1 address_4_reg_2_ ( .D(N131), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[2]) );
  DFFARX1 address_4_reg_1_ ( .D(N130), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[1]) );
  DFFARX1 address_4_reg_0_ ( .D(N129), .CLK(clk), .RSTB(rst_n), .Q(
        address_4[0]) );
  DFFARX1 address_2_reg_15_ ( .D(N176), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[15]) );
  DFFARX1 address_2_reg_14_ ( .D(N175), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[14]) );
  DFFARX1 address_2_reg_13_ ( .D(N174), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[13]) );
  DFFARX1 address_2_reg_12_ ( .D(N173), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[12]) );
  DFFARX1 address_2_reg_11_ ( .D(N172), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[11]) );
  DFFARX1 address_2_reg_10_ ( .D(N171), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[10]) );
  DFFARX1 address_2_reg_9_ ( .D(N170), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[9]) );
  DFFARX1 address_2_reg_8_ ( .D(N169), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[8]) );
  DFFARX1 address_2_reg_7_ ( .D(N168), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[7]) );
  DFFARX1 address_2_reg_6_ ( .D(N167), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[6]) );
  DFFARX1 address_2_reg_5_ ( .D(N166), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[5]) );
  DFFARX1 address_2_reg_4_ ( .D(N165), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[4]) );
  DFFARX1 address_2_reg_3_ ( .D(N164), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[3]) );
  DFFARX1 address_2_reg_2_ ( .D(N163), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[2]) );
  DFFARX1 address_2_reg_1_ ( .D(N162), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[1]) );
  DFFARX1 address_2_reg_0_ ( .D(N161), .CLK(clk), .RSTB(rst_n), .Q(
        address_2[0]) );
  DFFARX1 write_read_3_reg ( .D(N725), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_3) );
  DFFARX1 write_read_4_reg ( .D(N724), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_4) );
  DFFARX1 write_read_5_reg ( .D(N723), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_5) );
  DFFARX1 write_read_6_reg ( .D(N722), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_6) );
  DFFARX1 write_read_7_reg ( .D(N721), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_7) );
  DFFARX1 address_0_reg_15_ ( .D(N208), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[15]) );
  DFFARX1 address_0_reg_14_ ( .D(N207), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[14]) );
  DFFARX1 address_0_reg_13_ ( .D(N206), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[13]) );
  DFFARX1 address_0_reg_12_ ( .D(N205), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[12]) );
  DFFARX1 address_0_reg_11_ ( .D(N204), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[11]) );
  DFFARX1 address_0_reg_10_ ( .D(N203), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[10]) );
  DFFARX1 address_0_reg_9_ ( .D(N202), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[9]) );
  DFFARX1 address_0_reg_8_ ( .D(N201), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[8]) );
  DFFARX1 address_0_reg_7_ ( .D(N200), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[7]) );
  DFFARX1 address_0_reg_6_ ( .D(N199), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[6]) );
  DFFARX1 address_0_reg_5_ ( .D(N198), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[5]) );
  DFFARX1 address_0_reg_4_ ( .D(N197), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[4]) );
  DFFARX1 address_0_reg_3_ ( .D(N196), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[3]) );
  DFFARX1 address_0_reg_2_ ( .D(N195), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[2]) );
  DFFARX1 address_0_reg_1_ ( .D(N194), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[1]) );
  DFFARX1 address_0_reg_0_ ( .D(N193), .CLK(clk), .RSTB(rst_n), .Q(
        address_0[0]) );
  DFFARX1 address_1_reg_15_ ( .D(N192), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[15]) );
  DFFARX1 address_1_reg_14_ ( .D(N191), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[14]) );
  DFFARX1 address_1_reg_13_ ( .D(N190), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[13]) );
  DFFARX1 address_1_reg_12_ ( .D(N189), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[12]) );
  DFFARX1 address_1_reg_11_ ( .D(N188), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[11]) );
  DFFARX1 address_1_reg_10_ ( .D(N187), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[10]) );
  DFFARX1 address_1_reg_9_ ( .D(N186), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[9]) );
  DFFARX1 address_1_reg_8_ ( .D(N185), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[8]) );
  DFFARX1 address_1_reg_7_ ( .D(N184), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[7]) );
  DFFARX1 address_1_reg_6_ ( .D(N183), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[6]) );
  DFFARX1 address_1_reg_5_ ( .D(N182), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[5]) );
  DFFARX1 address_1_reg_4_ ( .D(N181), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[4]) );
  DFFARX1 address_1_reg_3_ ( .D(N180), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[3]) );
  DFFARX1 address_1_reg_2_ ( .D(N179), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[2]) );
  DFFARX1 address_1_reg_1_ ( .D(N178), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[1]) );
  DFFARX1 address_1_reg_0_ ( .D(N177), .CLK(clk), .RSTB(rst_n), .Q(
        address_1[0]) );
  DFFARX1 address_3_reg_15_ ( .D(N160), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[15]) );
  DFFARX1 address_3_reg_14_ ( .D(N159), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[14]) );
  DFFARX1 address_3_reg_13_ ( .D(N158), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[13]) );
  DFFARX1 address_3_reg_12_ ( .D(N157), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[12]) );
  DFFARX1 address_3_reg_11_ ( .D(N156), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[11]) );
  DFFARX1 address_3_reg_10_ ( .D(N155), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[10]) );
  DFFARX1 address_3_reg_9_ ( .D(N154), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[9]) );
  DFFARX1 address_3_reg_8_ ( .D(N153), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[8]) );
  DFFARX1 address_3_reg_7_ ( .D(N152), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[7]) );
  DFFARX1 address_3_reg_6_ ( .D(N151), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[6]) );
  DFFARX1 address_3_reg_5_ ( .D(N150), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[5]) );
  DFFARX1 address_3_reg_4_ ( .D(N149), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[4]) );
  DFFARX1 address_3_reg_3_ ( .D(N148), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[3]) );
  DFFARX1 address_3_reg_2_ ( .D(N147), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[2]) );
  DFFARX1 address_3_reg_1_ ( .D(N146), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[1]) );
  DFFARX1 address_3_reg_0_ ( .D(N145), .CLK(clk), .RSTB(rst_n), .Q(
        address_3[0]) );
  DFFARX1 write_read_1_reg ( .D(N727), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_1) );
  DFFARX1 write_read_2_reg ( .D(N726), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_2) );
  DFFARX1 write_read_0_reg ( .D(N728), .CLK(clk), .RSTB(rst_n), .Q(
        write_read_0) );
  DFFARX1 rdata_mbist_reg_63_ ( .D(N79), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[63]) );
  DFFARX1 rdata_mbist_reg_62_ ( .D(N78), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[62]) );
  DFFARX1 rdata_mbist_reg_61_ ( .D(N77), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[61]) );
  DFFARX1 rdata_mbist_reg_60_ ( .D(N76), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[60]) );
  DFFARX1 rdata_mbist_reg_59_ ( .D(N75), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[59]) );
  DFFARX1 rdata_mbist_reg_58_ ( .D(N74), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[58]) );
  DFFARX1 rdata_mbist_reg_57_ ( .D(N73), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[57]) );
  DFFARX1 rdata_mbist_reg_56_ ( .D(N72), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[56]) );
  DFFARX1 rdata_mbist_reg_55_ ( .D(N71), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[55]) );
  DFFARX1 rdata_mbist_reg_54_ ( .D(N70), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[54]) );
  DFFARX1 rdata_mbist_reg_53_ ( .D(N69), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[53]) );
  DFFARX1 rdata_mbist_reg_52_ ( .D(N68), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[52]) );
  DFFARX1 rdata_mbist_reg_51_ ( .D(N67), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[51]) );
  DFFARX1 rdata_mbist_reg_50_ ( .D(N66), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[50]) );
  DFFARX1 rdata_mbist_reg_49_ ( .D(N65), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[49]) );
  DFFARX1 rdata_mbist_reg_48_ ( .D(N64), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[48]) );
  DFFARX1 rdata_mbist_reg_47_ ( .D(N63), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[47]) );
  DFFARX1 rdata_mbist_reg_46_ ( .D(N62), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[46]) );
  DFFARX1 rdata_mbist_reg_45_ ( .D(N61), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[45]) );
  DFFARX1 rdata_mbist_reg_44_ ( .D(N60), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[44]) );
  DFFARX1 rdata_mbist_reg_43_ ( .D(N59), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[43]) );
  DFFARX1 rdata_mbist_reg_42_ ( .D(N58), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[42]) );
  DFFARX1 rdata_mbist_reg_41_ ( .D(N57), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[41]) );
  DFFARX1 rdata_mbist_reg_40_ ( .D(N56), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[40]) );
  DFFARX1 rdata_mbist_reg_39_ ( .D(N55), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[39]) );
  DFFARX1 rdata_mbist_reg_38_ ( .D(N54), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[38]) );
  DFFARX1 rdata_mbist_reg_37_ ( .D(N53), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[37]) );
  DFFARX1 rdata_mbist_reg_36_ ( .D(N52), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[36]) );
  DFFARX1 rdata_mbist_reg_35_ ( .D(N51), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[35]) );
  DFFARX1 rdata_mbist_reg_34_ ( .D(N50), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[34]) );
  DFFARX1 rdata_mbist_reg_33_ ( .D(N49), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[33]) );
  DFFARX1 rdata_mbist_reg_32_ ( .D(N48), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[32]) );
  DFFARX1 rdata_mbist_reg_31_ ( .D(N47), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[31]) );
  DFFARX1 rdata_mbist_reg_30_ ( .D(N46), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[30]) );
  DFFARX1 rdata_mbist_reg_29_ ( .D(N45), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[29]) );
  DFFARX1 rdata_mbist_reg_28_ ( .D(N44), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[28]) );
  DFFARX1 rdata_mbist_reg_27_ ( .D(N43), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[27]) );
  DFFARX1 rdata_mbist_reg_26_ ( .D(N42), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[26]) );
  DFFARX1 rdata_mbist_reg_25_ ( .D(N41), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[25]) );
  DFFARX1 rdata_mbist_reg_24_ ( .D(N40), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[24]) );
  DFFARX1 rdata_mbist_reg_23_ ( .D(N39), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[23]) );
  DFFARX1 rdata_mbist_reg_22_ ( .D(N38), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[22]) );
  DFFARX1 rdata_mbist_reg_21_ ( .D(N37), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[21]) );
  DFFARX1 rdata_mbist_reg_20_ ( .D(N36), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[20]) );
  DFFARX1 rdata_mbist_reg_19_ ( .D(N35), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[19]) );
  DFFARX1 rdata_mbist_reg_18_ ( .D(N34), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[18]) );
  DFFARX1 rdata_mbist_reg_17_ ( .D(N33), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[17]) );
  DFFARX1 rdata_mbist_reg_16_ ( .D(N32), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[16]) );
  DFFARX1 rdata_mbist_reg_15_ ( .D(N31), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[15]) );
  DFFARX1 rdata_mbist_reg_14_ ( .D(N30), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[14]) );
  DFFARX1 rdata_mbist_reg_13_ ( .D(N29), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[13]) );
  DFFARX1 rdata_mbist_reg_12_ ( .D(N28), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[12]) );
  DFFARX1 rdata_mbist_reg_11_ ( .D(N27), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[11]) );
  DFFARX1 rdata_mbist_reg_10_ ( .D(N26), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[10]) );
  DFFARX1 rdata_mbist_reg_9_ ( .D(N25), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[9]) );
  DFFARX1 rdata_mbist_reg_8_ ( .D(N24), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[8]) );
  DFFARX1 rdata_mbist_reg_7_ ( .D(N23), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[7]) );
  DFFARX1 rdata_mbist_reg_6_ ( .D(N22), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[6]) );
  DFFARX1 rdata_mbist_reg_5_ ( .D(N21), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[5]) );
  DFFARX1 rdata_mbist_reg_4_ ( .D(N20), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[4]) );
  DFFARX1 rdata_mbist_reg_3_ ( .D(N19), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[3]) );
  DFFARX1 rdata_mbist_reg_2_ ( .D(N18), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[2]) );
  DFFARX1 rdata_mbist_reg_1_ ( .D(N17), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[1]) );
  DFFARX1 rdata_mbist_reg_0_ ( .D(N16), .CLK(clk), .RSTB(rst_n), .Q(
        rdata_mbist[0]) );
  DFFARX1 wdata_7_reg_63_ ( .D(N272), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[63])
         );
  DFFARX1 wdata_7_reg_62_ ( .D(N271), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[62])
         );
  DFFARX1 wdata_7_reg_61_ ( .D(N270), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[61])
         );
  DFFARX1 wdata_7_reg_60_ ( .D(N269), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[60])
         );
  DFFARX1 wdata_7_reg_59_ ( .D(N268), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[59])
         );
  DFFARX1 wdata_7_reg_58_ ( .D(N267), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[58])
         );
  DFFARX1 wdata_7_reg_57_ ( .D(N266), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[57])
         );
  DFFARX1 wdata_7_reg_56_ ( .D(N265), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[56])
         );
  DFFARX1 wdata_7_reg_55_ ( .D(N264), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[55])
         );
  DFFARX1 wdata_7_reg_54_ ( .D(N263), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[54])
         );
  DFFARX1 wdata_7_reg_53_ ( .D(N262), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[53])
         );
  DFFARX1 wdata_7_reg_52_ ( .D(N261), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[52])
         );
  DFFARX1 wdata_7_reg_51_ ( .D(N260), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[51])
         );
  DFFARX1 wdata_7_reg_50_ ( .D(N259), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[50])
         );
  DFFARX1 wdata_7_reg_49_ ( .D(N258), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[49])
         );
  DFFARX1 wdata_7_reg_48_ ( .D(N257), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[48])
         );
  DFFARX1 wdata_7_reg_47_ ( .D(N256), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[47])
         );
  DFFARX1 wdata_7_reg_46_ ( .D(N255), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[46])
         );
  DFFARX1 wdata_7_reg_45_ ( .D(N254), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[45])
         );
  DFFARX1 wdata_7_reg_44_ ( .D(N253), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[44])
         );
  DFFARX1 wdata_7_reg_43_ ( .D(N252), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[43])
         );
  DFFARX1 wdata_7_reg_42_ ( .D(N251), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[42])
         );
  DFFARX1 wdata_7_reg_41_ ( .D(N250), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[41])
         );
  DFFARX1 wdata_7_reg_40_ ( .D(N249), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[40])
         );
  DFFARX1 wdata_7_reg_39_ ( .D(N248), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[39])
         );
  DFFARX1 wdata_7_reg_38_ ( .D(N247), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[38])
         );
  DFFARX1 wdata_7_reg_37_ ( .D(N246), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[37])
         );
  DFFARX1 wdata_7_reg_36_ ( .D(N245), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[36])
         );
  DFFARX1 wdata_7_reg_35_ ( .D(N244), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[35])
         );
  DFFARX1 wdata_7_reg_34_ ( .D(N243), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[34])
         );
  DFFARX1 wdata_7_reg_33_ ( .D(N242), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[33])
         );
  DFFARX1 wdata_7_reg_32_ ( .D(N241), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[32])
         );
  DFFARX1 wdata_7_reg_31_ ( .D(N240), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[31])
         );
  DFFARX1 wdata_7_reg_30_ ( .D(N239), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[30])
         );
  DFFARX1 wdata_7_reg_29_ ( .D(N238), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[29])
         );
  DFFARX1 wdata_7_reg_28_ ( .D(N237), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[28])
         );
  DFFARX1 wdata_7_reg_27_ ( .D(N236), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[27])
         );
  DFFARX1 wdata_7_reg_26_ ( .D(N235), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[26])
         );
  DFFARX1 wdata_7_reg_25_ ( .D(N234), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[25])
         );
  DFFARX1 wdata_7_reg_24_ ( .D(N233), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[24])
         );
  DFFARX1 wdata_7_reg_23_ ( .D(N232), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[23])
         );
  DFFARX1 wdata_7_reg_22_ ( .D(N231), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[22])
         );
  DFFARX1 wdata_7_reg_21_ ( .D(N230), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[21])
         );
  DFFARX1 wdata_7_reg_20_ ( .D(N229), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[20])
         );
  DFFARX1 wdata_7_reg_19_ ( .D(N228), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[19])
         );
  DFFARX1 wdata_7_reg_18_ ( .D(N227), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[18])
         );
  DFFARX1 wdata_7_reg_17_ ( .D(N226), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[17])
         );
  DFFARX1 wdata_7_reg_16_ ( .D(N225), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[16])
         );
  DFFARX1 wdata_7_reg_15_ ( .D(N224), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[15])
         );
  DFFARX1 wdata_7_reg_14_ ( .D(N223), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[14])
         );
  DFFARX1 wdata_7_reg_13_ ( .D(N222), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[13])
         );
  DFFARX1 wdata_7_reg_12_ ( .D(N221), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[12])
         );
  DFFARX1 wdata_7_reg_11_ ( .D(N220), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[11])
         );
  DFFARX1 wdata_7_reg_10_ ( .D(N219), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[10])
         );
  DFFARX1 wdata_7_reg_9_ ( .D(N218), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[9])
         );
  DFFARX1 wdata_7_reg_8_ ( .D(N217), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[8])
         );
  DFFARX1 wdata_7_reg_7_ ( .D(N216), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[7])
         );
  DFFARX1 wdata_7_reg_6_ ( .D(N215), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[6])
         );
  DFFARX1 wdata_7_reg_5_ ( .D(N214), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[5])
         );
  DFFARX1 wdata_7_reg_4_ ( .D(N213), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[4])
         );
  DFFARX1 wdata_7_reg_3_ ( .D(N212), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[3])
         );
  DFFARX1 wdata_7_reg_2_ ( .D(N211), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[2])
         );
  DFFARX1 wdata_7_reg_1_ ( .D(N210), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[1])
         );
  DFFARX1 wdata_7_reg_0_ ( .D(N209), .CLK(clk), .RSTB(rst_n), .Q(wdata_7[0])
         );
  DFFARX1 wdata_6_reg_63_ ( .D(N336), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[63])
         );
  DFFARX1 wdata_6_reg_62_ ( .D(N335), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[62])
         );
  DFFARX1 wdata_6_reg_61_ ( .D(N334), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[61])
         );
  DFFARX1 wdata_6_reg_60_ ( .D(N333), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[60])
         );
  DFFARX1 wdata_6_reg_59_ ( .D(N332), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[59])
         );
  DFFARX1 wdata_6_reg_58_ ( .D(N331), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[58])
         );
  DFFARX1 wdata_6_reg_57_ ( .D(N330), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[57])
         );
  DFFARX1 wdata_6_reg_56_ ( .D(N329), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[56])
         );
  DFFARX1 wdata_6_reg_55_ ( .D(N328), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[55])
         );
  DFFARX1 wdata_6_reg_54_ ( .D(N327), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[54])
         );
  DFFARX1 wdata_6_reg_53_ ( .D(N326), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[53])
         );
  DFFARX1 wdata_6_reg_52_ ( .D(N325), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[52])
         );
  DFFARX1 wdata_6_reg_51_ ( .D(N324), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[51])
         );
  DFFARX1 wdata_6_reg_50_ ( .D(N323), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[50])
         );
  DFFARX1 wdata_6_reg_49_ ( .D(N322), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[49])
         );
  DFFARX1 wdata_6_reg_48_ ( .D(N321), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[48])
         );
  DFFARX1 wdata_6_reg_47_ ( .D(N320), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[47])
         );
  DFFARX1 wdata_6_reg_46_ ( .D(N319), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[46])
         );
  DFFARX1 wdata_6_reg_45_ ( .D(N318), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[45])
         );
  DFFARX1 wdata_6_reg_44_ ( .D(N317), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[44])
         );
  DFFARX1 wdata_6_reg_43_ ( .D(N316), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[43])
         );
  DFFARX1 wdata_6_reg_42_ ( .D(N315), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[42])
         );
  DFFARX1 wdata_6_reg_41_ ( .D(N314), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[41])
         );
  DFFARX1 wdata_6_reg_40_ ( .D(N313), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[40])
         );
  DFFARX1 wdata_6_reg_39_ ( .D(N312), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[39])
         );
  DFFARX1 wdata_6_reg_38_ ( .D(N311), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[38])
         );
  DFFARX1 wdata_6_reg_37_ ( .D(N310), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[37])
         );
  DFFARX1 wdata_6_reg_36_ ( .D(N309), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[36])
         );
  DFFARX1 wdata_6_reg_35_ ( .D(N308), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[35])
         );
  DFFARX1 wdata_6_reg_34_ ( .D(N307), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[34])
         );
  DFFARX1 wdata_6_reg_33_ ( .D(N306), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[33])
         );
  DFFARX1 wdata_6_reg_32_ ( .D(N305), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[32])
         );
  DFFARX1 wdata_6_reg_31_ ( .D(N304), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[31])
         );
  DFFARX1 wdata_6_reg_30_ ( .D(N303), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[30])
         );
  DFFARX1 wdata_6_reg_29_ ( .D(N302), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[29])
         );
  DFFARX1 wdata_6_reg_28_ ( .D(N301), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[28])
         );
  DFFARX1 wdata_6_reg_27_ ( .D(N300), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[27])
         );
  DFFARX1 wdata_6_reg_26_ ( .D(N299), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[26])
         );
  DFFARX1 wdata_6_reg_25_ ( .D(N298), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[25])
         );
  DFFARX1 wdata_6_reg_24_ ( .D(N297), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[24])
         );
  DFFARX1 wdata_6_reg_23_ ( .D(N296), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[23])
         );
  DFFARX1 wdata_6_reg_22_ ( .D(N295), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[22])
         );
  DFFARX1 wdata_6_reg_21_ ( .D(N294), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[21])
         );
  DFFARX1 wdata_6_reg_20_ ( .D(N293), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[20])
         );
  DFFARX1 wdata_6_reg_19_ ( .D(N292), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[19])
         );
  DFFARX1 wdata_6_reg_18_ ( .D(N291), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[18])
         );
  DFFARX1 wdata_6_reg_17_ ( .D(N290), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[17])
         );
  DFFARX1 wdata_6_reg_16_ ( .D(N289), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[16])
         );
  DFFARX1 wdata_6_reg_15_ ( .D(N288), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[15])
         );
  DFFARX1 wdata_6_reg_14_ ( .D(N287), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[14])
         );
  DFFARX1 wdata_6_reg_13_ ( .D(N286), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[13])
         );
  DFFARX1 wdata_6_reg_12_ ( .D(N285), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[12])
         );
  DFFARX1 wdata_6_reg_11_ ( .D(N284), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[11])
         );
  DFFARX1 wdata_6_reg_10_ ( .D(N283), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[10])
         );
  DFFARX1 wdata_6_reg_9_ ( .D(N282), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[9])
         );
  DFFARX1 wdata_6_reg_8_ ( .D(N281), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[8])
         );
  DFFARX1 wdata_6_reg_7_ ( .D(N280), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[7])
         );
  DFFARX1 wdata_6_reg_6_ ( .D(N279), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[6])
         );
  DFFARX1 wdata_6_reg_5_ ( .D(N278), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[5])
         );
  DFFARX1 wdata_6_reg_4_ ( .D(N277), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[4])
         );
  DFFARX1 wdata_6_reg_3_ ( .D(N276), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[3])
         );
  DFFARX1 wdata_6_reg_2_ ( .D(N275), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[2])
         );
  DFFARX1 wdata_6_reg_1_ ( .D(N274), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[1])
         );
  DFFARX1 wdata_6_reg_0_ ( .D(N273), .CLK(clk), .RSTB(rst_n), .Q(wdata_6[0])
         );
  DFFARX1 wdata_5_reg_63_ ( .D(N400), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[63])
         );
  DFFARX1 wdata_5_reg_62_ ( .D(N399), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[62])
         );
  DFFARX1 wdata_5_reg_61_ ( .D(N398), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[61])
         );
  DFFARX1 wdata_5_reg_60_ ( .D(N397), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[60])
         );
  DFFARX1 wdata_5_reg_59_ ( .D(N396), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[59])
         );
  DFFARX1 wdata_5_reg_58_ ( .D(N395), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[58])
         );
  DFFARX1 wdata_5_reg_57_ ( .D(N394), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[57])
         );
  DFFARX1 wdata_5_reg_56_ ( .D(N393), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[56])
         );
  DFFARX1 wdata_5_reg_55_ ( .D(N392), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[55])
         );
  DFFARX1 wdata_5_reg_54_ ( .D(N391), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[54])
         );
  DFFARX1 wdata_5_reg_53_ ( .D(N390), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[53])
         );
  DFFARX1 wdata_5_reg_52_ ( .D(N389), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[52])
         );
  DFFARX1 wdata_5_reg_51_ ( .D(N388), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[51])
         );
  DFFARX1 wdata_5_reg_50_ ( .D(N387), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[50])
         );
  DFFARX1 wdata_5_reg_49_ ( .D(N386), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[49])
         );
  DFFARX1 wdata_5_reg_48_ ( .D(N385), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[48])
         );
  DFFARX1 wdata_5_reg_47_ ( .D(N384), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[47])
         );
  DFFARX1 wdata_5_reg_46_ ( .D(N383), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[46])
         );
  DFFARX1 wdata_5_reg_45_ ( .D(N382), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[45])
         );
  DFFARX1 wdata_5_reg_44_ ( .D(N381), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[44])
         );
  DFFARX1 wdata_5_reg_43_ ( .D(N380), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[43])
         );
  DFFARX1 wdata_5_reg_42_ ( .D(N379), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[42])
         );
  DFFARX1 wdata_5_reg_41_ ( .D(N378), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[41])
         );
  DFFARX1 wdata_5_reg_40_ ( .D(N377), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[40])
         );
  DFFARX1 wdata_5_reg_39_ ( .D(N376), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[39])
         );
  DFFARX1 wdata_5_reg_38_ ( .D(N375), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[38])
         );
  DFFARX1 wdata_5_reg_37_ ( .D(N374), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[37])
         );
  DFFARX1 wdata_5_reg_36_ ( .D(N373), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[36])
         );
  DFFARX1 wdata_5_reg_35_ ( .D(N372), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[35])
         );
  DFFARX1 wdata_5_reg_34_ ( .D(N371), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[34])
         );
  DFFARX1 wdata_5_reg_33_ ( .D(N370), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[33])
         );
  DFFARX1 wdata_5_reg_32_ ( .D(N369), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[32])
         );
  DFFARX1 wdata_5_reg_31_ ( .D(N368), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[31])
         );
  DFFARX1 wdata_5_reg_30_ ( .D(N367), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[30])
         );
  DFFARX1 wdata_5_reg_29_ ( .D(N366), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[29])
         );
  DFFARX1 wdata_5_reg_28_ ( .D(N365), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[28])
         );
  DFFARX1 wdata_5_reg_27_ ( .D(N364), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[27])
         );
  DFFARX1 wdata_5_reg_26_ ( .D(N363), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[26])
         );
  DFFARX1 wdata_5_reg_25_ ( .D(N362), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[25])
         );
  DFFARX1 wdata_5_reg_24_ ( .D(N361), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[24])
         );
  DFFARX1 wdata_5_reg_23_ ( .D(N360), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[23])
         );
  DFFARX1 wdata_5_reg_22_ ( .D(N359), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[22])
         );
  DFFARX1 wdata_5_reg_21_ ( .D(N358), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[21])
         );
  DFFARX1 wdata_5_reg_20_ ( .D(N357), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[20])
         );
  DFFARX1 wdata_5_reg_19_ ( .D(N356), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[19])
         );
  DFFARX1 wdata_5_reg_18_ ( .D(N355), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[18])
         );
  DFFARX1 wdata_5_reg_17_ ( .D(N354), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[17])
         );
  DFFARX1 wdata_5_reg_16_ ( .D(N353), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[16])
         );
  DFFARX1 wdata_5_reg_15_ ( .D(N352), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[15])
         );
  DFFARX1 wdata_5_reg_14_ ( .D(N351), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[14])
         );
  DFFARX1 wdata_5_reg_13_ ( .D(N350), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[13])
         );
  DFFARX1 wdata_5_reg_12_ ( .D(N349), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[12])
         );
  DFFARX1 wdata_5_reg_11_ ( .D(N348), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[11])
         );
  DFFARX1 wdata_5_reg_10_ ( .D(N347), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[10])
         );
  DFFARX1 wdata_5_reg_9_ ( .D(N346), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[9])
         );
  DFFARX1 wdata_5_reg_8_ ( .D(N345), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[8])
         );
  DFFARX1 wdata_5_reg_7_ ( .D(N344), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[7])
         );
  DFFARX1 wdata_5_reg_6_ ( .D(N343), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[6])
         );
  DFFARX1 wdata_5_reg_5_ ( .D(N342), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[5])
         );
  DFFARX1 wdata_5_reg_4_ ( .D(N341), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[4])
         );
  DFFARX1 wdata_5_reg_3_ ( .D(N340), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[3])
         );
  DFFARX1 wdata_5_reg_2_ ( .D(N339), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[2])
         );
  DFFARX1 wdata_5_reg_1_ ( .D(N338), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[1])
         );
  DFFARX1 wdata_5_reg_0_ ( .D(N337), .CLK(clk), .RSTB(rst_n), .Q(wdata_5[0])
         );
  DFFARX1 wdata_4_reg_63_ ( .D(N464), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[63])
         );
  DFFARX1 wdata_4_reg_62_ ( .D(N463), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[62])
         );
  DFFARX1 wdata_4_reg_61_ ( .D(N462), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[61])
         );
  DFFARX1 wdata_4_reg_60_ ( .D(N461), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[60])
         );
  DFFARX1 wdata_4_reg_59_ ( .D(N460), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[59])
         );
  DFFARX1 wdata_4_reg_58_ ( .D(N459), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[58])
         );
  DFFARX1 wdata_4_reg_57_ ( .D(N458), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[57])
         );
  DFFARX1 wdata_4_reg_56_ ( .D(N457), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[56])
         );
  DFFARX1 wdata_4_reg_55_ ( .D(N456), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[55])
         );
  DFFARX1 wdata_4_reg_54_ ( .D(N455), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[54])
         );
  DFFARX1 wdata_4_reg_53_ ( .D(N454), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[53])
         );
  DFFARX1 wdata_4_reg_52_ ( .D(N453), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[52])
         );
  DFFARX1 wdata_4_reg_51_ ( .D(N452), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[51])
         );
  DFFARX1 wdata_4_reg_50_ ( .D(N451), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[50])
         );
  DFFARX1 wdata_4_reg_49_ ( .D(N450), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[49])
         );
  DFFARX1 wdata_4_reg_48_ ( .D(N449), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[48])
         );
  DFFARX1 wdata_4_reg_47_ ( .D(N448), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[47])
         );
  DFFARX1 wdata_4_reg_46_ ( .D(N447), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[46])
         );
  DFFARX1 wdata_4_reg_45_ ( .D(N446), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[45])
         );
  DFFARX1 wdata_4_reg_44_ ( .D(N445), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[44])
         );
  DFFARX1 wdata_4_reg_43_ ( .D(N444), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[43])
         );
  DFFARX1 wdata_4_reg_42_ ( .D(N443), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[42])
         );
  DFFARX1 wdata_4_reg_41_ ( .D(N442), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[41])
         );
  DFFARX1 wdata_4_reg_40_ ( .D(N441), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[40])
         );
  DFFARX1 wdata_4_reg_39_ ( .D(N440), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[39])
         );
  DFFARX1 wdata_4_reg_38_ ( .D(N439), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[38])
         );
  DFFARX1 wdata_4_reg_37_ ( .D(N438), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[37])
         );
  DFFARX1 wdata_4_reg_36_ ( .D(N437), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[36])
         );
  DFFARX1 wdata_4_reg_35_ ( .D(N436), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[35])
         );
  DFFARX1 wdata_4_reg_34_ ( .D(N435), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[34])
         );
  DFFARX1 wdata_4_reg_33_ ( .D(N434), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[33])
         );
  DFFARX1 wdata_4_reg_32_ ( .D(N433), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[32])
         );
  DFFARX1 wdata_4_reg_31_ ( .D(N432), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[31])
         );
  DFFARX1 wdata_4_reg_30_ ( .D(N431), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[30])
         );
  DFFARX1 wdata_4_reg_29_ ( .D(N430), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[29])
         );
  DFFARX1 wdata_4_reg_28_ ( .D(N429), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[28])
         );
  DFFARX1 wdata_4_reg_27_ ( .D(N428), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[27])
         );
  DFFARX1 wdata_4_reg_26_ ( .D(N427), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[26])
         );
  DFFARX1 wdata_4_reg_25_ ( .D(N426), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[25])
         );
  DFFARX1 wdata_4_reg_24_ ( .D(N425), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[24])
         );
  DFFARX1 wdata_4_reg_23_ ( .D(N424), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[23])
         );
  DFFARX1 wdata_4_reg_22_ ( .D(N423), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[22])
         );
  DFFARX1 wdata_4_reg_21_ ( .D(N422), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[21])
         );
  DFFARX1 wdata_4_reg_20_ ( .D(N421), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[20])
         );
  DFFARX1 wdata_4_reg_19_ ( .D(N420), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[19])
         );
  DFFARX1 wdata_4_reg_18_ ( .D(N419), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[18])
         );
  DFFARX1 wdata_4_reg_17_ ( .D(N418), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[17])
         );
  DFFARX1 wdata_4_reg_16_ ( .D(N417), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[16])
         );
  DFFARX1 wdata_4_reg_15_ ( .D(N416), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[15])
         );
  DFFARX1 wdata_4_reg_14_ ( .D(N415), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[14])
         );
  DFFARX1 wdata_4_reg_13_ ( .D(N414), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[13])
         );
  DFFARX1 wdata_4_reg_12_ ( .D(N413), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[12])
         );
  DFFARX1 wdata_4_reg_11_ ( .D(N412), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[11])
         );
  DFFARX1 wdata_4_reg_10_ ( .D(N411), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[10])
         );
  DFFARX1 wdata_4_reg_9_ ( .D(N410), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[9])
         );
  DFFARX1 wdata_4_reg_8_ ( .D(N409), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[8])
         );
  DFFARX1 wdata_4_reg_7_ ( .D(N408), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[7])
         );
  DFFARX1 wdata_4_reg_6_ ( .D(N407), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[6])
         );
  DFFARX1 wdata_4_reg_5_ ( .D(N406), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[5])
         );
  DFFARX1 wdata_4_reg_4_ ( .D(N405), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[4])
         );
  DFFARX1 wdata_4_reg_3_ ( .D(N404), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[3])
         );
  DFFARX1 wdata_4_reg_2_ ( .D(N403), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[2])
         );
  DFFARX1 wdata_4_reg_1_ ( .D(N402), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[1])
         );
  DFFARX1 wdata_4_reg_0_ ( .D(N401), .CLK(clk), .RSTB(rst_n), .Q(wdata_4[0])
         );
  DFFARX1 wdata_3_reg_63_ ( .D(N528), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[63])
         );
  DFFARX1 wdata_3_reg_62_ ( .D(N527), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[62])
         );
  DFFARX1 wdata_3_reg_61_ ( .D(N526), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[61])
         );
  DFFARX1 wdata_3_reg_60_ ( .D(N525), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[60])
         );
  DFFARX1 wdata_3_reg_59_ ( .D(N524), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[59])
         );
  DFFARX1 wdata_3_reg_58_ ( .D(N523), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[58])
         );
  DFFARX1 wdata_3_reg_57_ ( .D(N522), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[57])
         );
  DFFARX1 wdata_3_reg_56_ ( .D(N521), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[56])
         );
  DFFARX1 wdata_3_reg_55_ ( .D(N520), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[55])
         );
  DFFARX1 wdata_3_reg_54_ ( .D(N519), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[54])
         );
  DFFARX1 wdata_3_reg_53_ ( .D(N518), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[53])
         );
  DFFARX1 wdata_3_reg_52_ ( .D(N517), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[52])
         );
  DFFARX1 wdata_3_reg_51_ ( .D(N516), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[51])
         );
  DFFARX1 wdata_3_reg_50_ ( .D(N515), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[50])
         );
  DFFARX1 wdata_3_reg_49_ ( .D(N514), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[49])
         );
  DFFARX1 wdata_3_reg_48_ ( .D(N513), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[48])
         );
  DFFARX1 wdata_3_reg_47_ ( .D(N512), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[47])
         );
  DFFARX1 wdata_3_reg_46_ ( .D(N511), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[46])
         );
  DFFARX1 wdata_3_reg_45_ ( .D(N510), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[45])
         );
  DFFARX1 wdata_3_reg_44_ ( .D(N509), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[44])
         );
  DFFARX1 wdata_3_reg_43_ ( .D(N508), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[43])
         );
  DFFARX1 wdata_3_reg_42_ ( .D(N507), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[42])
         );
  DFFARX1 wdata_3_reg_41_ ( .D(N506), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[41])
         );
  DFFARX1 wdata_3_reg_40_ ( .D(N505), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[40])
         );
  DFFARX1 wdata_3_reg_39_ ( .D(N504), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[39])
         );
  DFFARX1 wdata_3_reg_38_ ( .D(N503), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[38])
         );
  DFFARX1 wdata_3_reg_37_ ( .D(N502), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[37])
         );
  DFFARX1 wdata_3_reg_36_ ( .D(N501), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[36])
         );
  DFFARX1 wdata_3_reg_35_ ( .D(N500), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[35])
         );
  DFFARX1 wdata_3_reg_34_ ( .D(N499), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[34])
         );
  DFFARX1 wdata_3_reg_33_ ( .D(N498), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[33])
         );
  DFFARX1 wdata_3_reg_32_ ( .D(N497), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[32])
         );
  DFFARX1 wdata_3_reg_31_ ( .D(N496), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[31])
         );
  DFFARX1 wdata_3_reg_30_ ( .D(N495), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[30])
         );
  DFFARX1 wdata_3_reg_29_ ( .D(N494), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[29])
         );
  DFFARX1 wdata_3_reg_28_ ( .D(N493), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[28])
         );
  DFFARX1 wdata_3_reg_27_ ( .D(N492), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[27])
         );
  DFFARX1 wdata_3_reg_26_ ( .D(N491), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[26])
         );
  DFFARX1 wdata_3_reg_25_ ( .D(N490), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[25])
         );
  DFFARX1 wdata_3_reg_24_ ( .D(N489), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[24])
         );
  DFFARX1 wdata_3_reg_23_ ( .D(N488), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[23])
         );
  DFFARX1 wdata_3_reg_22_ ( .D(N487), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[22])
         );
  DFFARX1 wdata_3_reg_21_ ( .D(N486), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[21])
         );
  DFFARX1 wdata_3_reg_20_ ( .D(N485), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[20])
         );
  DFFARX1 wdata_3_reg_19_ ( .D(N484), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[19])
         );
  DFFARX1 wdata_3_reg_18_ ( .D(N483), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[18])
         );
  DFFARX1 wdata_3_reg_17_ ( .D(N482), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[17])
         );
  DFFARX1 wdata_3_reg_16_ ( .D(N481), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[16])
         );
  DFFARX1 wdata_3_reg_15_ ( .D(N480), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[15])
         );
  DFFARX1 wdata_3_reg_14_ ( .D(N479), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[14])
         );
  DFFARX1 wdata_3_reg_13_ ( .D(N478), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[13])
         );
  DFFARX1 wdata_3_reg_12_ ( .D(N477), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[12])
         );
  DFFARX1 wdata_3_reg_11_ ( .D(N476), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[11])
         );
  DFFARX1 wdata_3_reg_10_ ( .D(N475), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[10])
         );
  DFFARX1 wdata_3_reg_9_ ( .D(N474), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[9])
         );
  DFFARX1 wdata_3_reg_8_ ( .D(N473), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[8])
         );
  DFFARX1 wdata_3_reg_7_ ( .D(N472), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[7])
         );
  DFFARX1 wdata_3_reg_6_ ( .D(N471), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[6])
         );
  DFFARX1 wdata_3_reg_5_ ( .D(N470), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[5])
         );
  DFFARX1 wdata_3_reg_4_ ( .D(N469), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[4])
         );
  DFFARX1 wdata_3_reg_3_ ( .D(N468), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[3])
         );
  DFFARX1 wdata_3_reg_2_ ( .D(N467), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[2])
         );
  DFFARX1 wdata_3_reg_1_ ( .D(N466), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[1])
         );
  DFFARX1 wdata_3_reg_0_ ( .D(N465), .CLK(clk), .RSTB(rst_n), .Q(wdata_3[0])
         );
  DFFARX1 wdata_2_reg_63_ ( .D(N592), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[63])
         );
  DFFARX1 wdata_2_reg_62_ ( .D(N591), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[62])
         );
  DFFARX1 wdata_2_reg_61_ ( .D(N590), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[61])
         );
  DFFARX1 wdata_2_reg_60_ ( .D(N589), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[60])
         );
  DFFARX1 wdata_2_reg_59_ ( .D(N588), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[59])
         );
  DFFARX1 wdata_2_reg_58_ ( .D(N587), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[58])
         );
  DFFARX1 wdata_2_reg_57_ ( .D(N586), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[57])
         );
  DFFARX1 wdata_2_reg_56_ ( .D(N585), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[56])
         );
  DFFARX1 wdata_2_reg_55_ ( .D(N584), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[55])
         );
  DFFARX1 wdata_2_reg_54_ ( .D(N583), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[54])
         );
  DFFARX1 wdata_2_reg_53_ ( .D(N582), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[53])
         );
  DFFARX1 wdata_2_reg_52_ ( .D(N581), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[52])
         );
  DFFARX1 wdata_2_reg_51_ ( .D(N580), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[51])
         );
  DFFARX1 wdata_2_reg_50_ ( .D(N579), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[50])
         );
  DFFARX1 wdata_2_reg_49_ ( .D(N578), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[49])
         );
  DFFARX1 wdata_2_reg_48_ ( .D(N577), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[48])
         );
  DFFARX1 wdata_2_reg_47_ ( .D(N576), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[47])
         );
  DFFARX1 wdata_2_reg_46_ ( .D(N575), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[46])
         );
  DFFARX1 wdata_2_reg_45_ ( .D(N574), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[45])
         );
  DFFARX1 wdata_2_reg_44_ ( .D(N573), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[44])
         );
  DFFARX1 wdata_2_reg_43_ ( .D(N572), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[43])
         );
  DFFARX1 wdata_2_reg_42_ ( .D(N571), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[42])
         );
  DFFARX1 wdata_2_reg_41_ ( .D(N570), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[41])
         );
  DFFARX1 wdata_2_reg_40_ ( .D(N569), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[40])
         );
  DFFARX1 wdata_2_reg_39_ ( .D(N568), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[39])
         );
  DFFARX1 wdata_2_reg_38_ ( .D(N567), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[38])
         );
  DFFARX1 wdata_2_reg_37_ ( .D(N566), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[37])
         );
  DFFARX1 wdata_2_reg_36_ ( .D(N565), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[36])
         );
  DFFARX1 wdata_2_reg_35_ ( .D(N564), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[35])
         );
  DFFARX1 wdata_2_reg_34_ ( .D(N563), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[34])
         );
  DFFARX1 wdata_2_reg_33_ ( .D(N562), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[33])
         );
  DFFARX1 wdata_2_reg_32_ ( .D(N561), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[32])
         );
  DFFARX1 wdata_2_reg_31_ ( .D(N560), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[31])
         );
  DFFARX1 wdata_2_reg_30_ ( .D(N559), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[30])
         );
  DFFARX1 wdata_2_reg_29_ ( .D(N558), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[29])
         );
  DFFARX1 wdata_2_reg_28_ ( .D(N557), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[28])
         );
  DFFARX1 wdata_2_reg_27_ ( .D(N556), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[27])
         );
  DFFARX1 wdata_2_reg_26_ ( .D(N555), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[26])
         );
  DFFARX1 wdata_2_reg_25_ ( .D(N554), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[25])
         );
  DFFARX1 wdata_2_reg_24_ ( .D(N553), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[24])
         );
  DFFARX1 wdata_2_reg_23_ ( .D(N552), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[23])
         );
  DFFARX1 wdata_2_reg_22_ ( .D(N551), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[22])
         );
  DFFARX1 wdata_2_reg_21_ ( .D(N550), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[21])
         );
  DFFARX1 wdata_2_reg_20_ ( .D(N549), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[20])
         );
  DFFARX1 wdata_2_reg_19_ ( .D(N548), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[19])
         );
  DFFARX1 wdata_2_reg_18_ ( .D(N547), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[18])
         );
  DFFARX1 wdata_2_reg_17_ ( .D(N546), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[17])
         );
  DFFARX1 wdata_2_reg_16_ ( .D(N545), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[16])
         );
  DFFARX1 wdata_2_reg_15_ ( .D(N544), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[15])
         );
  DFFARX1 wdata_2_reg_14_ ( .D(N543), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[14])
         );
  DFFARX1 wdata_2_reg_13_ ( .D(N542), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[13])
         );
  DFFARX1 wdata_2_reg_12_ ( .D(N541), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[12])
         );
  DFFARX1 wdata_2_reg_11_ ( .D(N540), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[11])
         );
  DFFARX1 wdata_2_reg_10_ ( .D(N539), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[10])
         );
  DFFARX1 wdata_2_reg_9_ ( .D(N538), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[9])
         );
  DFFARX1 wdata_2_reg_8_ ( .D(N537), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[8])
         );
  DFFARX1 wdata_2_reg_7_ ( .D(N536), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[7])
         );
  DFFARX1 wdata_2_reg_6_ ( .D(N535), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[6])
         );
  DFFARX1 wdata_2_reg_5_ ( .D(N534), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[5])
         );
  DFFARX1 wdata_2_reg_4_ ( .D(N533), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[4])
         );
  DFFARX1 wdata_2_reg_3_ ( .D(N532), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[3])
         );
  DFFARX1 wdata_2_reg_2_ ( .D(N531), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[2])
         );
  DFFARX1 wdata_2_reg_1_ ( .D(N530), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[1])
         );
  DFFARX1 wdata_2_reg_0_ ( .D(N529), .CLK(clk), .RSTB(rst_n), .Q(wdata_2[0])
         );
  DFFARX1 wdata_1_reg_63_ ( .D(N656), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[63])
         );
  DFFARX1 wdata_1_reg_62_ ( .D(N655), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[62])
         );
  DFFARX1 wdata_1_reg_61_ ( .D(N654), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[61])
         );
  DFFARX1 wdata_1_reg_60_ ( .D(N653), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[60])
         );
  DFFARX1 wdata_1_reg_59_ ( .D(N652), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[59])
         );
  DFFARX1 wdata_1_reg_58_ ( .D(N651), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[58])
         );
  DFFARX1 wdata_1_reg_57_ ( .D(N650), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[57])
         );
  DFFARX1 wdata_1_reg_56_ ( .D(N649), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[56])
         );
  DFFARX1 wdata_1_reg_55_ ( .D(N648), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[55])
         );
  DFFARX1 wdata_1_reg_54_ ( .D(N647), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[54])
         );
  DFFARX1 wdata_1_reg_53_ ( .D(N646), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[53])
         );
  DFFARX1 wdata_1_reg_52_ ( .D(N645), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[52])
         );
  DFFARX1 wdata_1_reg_51_ ( .D(N644), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[51])
         );
  DFFARX1 wdata_1_reg_50_ ( .D(N643), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[50])
         );
  DFFARX1 wdata_1_reg_49_ ( .D(N642), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[49])
         );
  DFFARX1 wdata_1_reg_48_ ( .D(N641), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[48])
         );
  DFFARX1 wdata_1_reg_47_ ( .D(N640), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[47])
         );
  DFFARX1 wdata_1_reg_46_ ( .D(N639), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[46])
         );
  DFFARX1 wdata_1_reg_45_ ( .D(N638), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[45])
         );
  DFFARX1 wdata_1_reg_44_ ( .D(N637), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[44])
         );
  DFFARX1 wdata_1_reg_43_ ( .D(N636), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[43])
         );
  DFFARX1 wdata_1_reg_42_ ( .D(N635), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[42])
         );
  DFFARX1 wdata_1_reg_41_ ( .D(N634), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[41])
         );
  DFFARX1 wdata_1_reg_40_ ( .D(N633), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[40])
         );
  DFFARX1 wdata_1_reg_39_ ( .D(N632), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[39])
         );
  DFFARX1 wdata_1_reg_38_ ( .D(N631), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[38])
         );
  DFFARX1 wdata_1_reg_37_ ( .D(N630), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[37])
         );
  DFFARX1 wdata_1_reg_36_ ( .D(N629), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[36])
         );
  DFFARX1 wdata_1_reg_35_ ( .D(N628), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[35])
         );
  DFFARX1 wdata_1_reg_34_ ( .D(N627), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[34])
         );
  DFFARX1 wdata_1_reg_33_ ( .D(N626), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[33])
         );
  DFFARX1 wdata_1_reg_32_ ( .D(N625), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[32])
         );
  DFFARX1 wdata_1_reg_31_ ( .D(N624), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[31])
         );
  DFFARX1 wdata_1_reg_30_ ( .D(N623), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[30])
         );
  DFFARX1 wdata_1_reg_29_ ( .D(N622), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[29])
         );
  DFFARX1 wdata_1_reg_28_ ( .D(N621), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[28])
         );
  DFFARX1 wdata_1_reg_27_ ( .D(N620), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[27])
         );
  DFFARX1 wdata_1_reg_26_ ( .D(N619), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[26])
         );
  DFFARX1 wdata_1_reg_25_ ( .D(N618), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[25])
         );
  DFFARX1 wdata_1_reg_24_ ( .D(N617), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[24])
         );
  DFFARX1 wdata_1_reg_23_ ( .D(N616), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[23])
         );
  DFFARX1 wdata_1_reg_22_ ( .D(N615), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[22])
         );
  DFFARX1 wdata_1_reg_21_ ( .D(N614), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[21])
         );
  DFFARX1 wdata_1_reg_20_ ( .D(N613), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[20])
         );
  DFFARX1 wdata_1_reg_19_ ( .D(N612), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[19])
         );
  DFFARX1 wdata_1_reg_18_ ( .D(N611), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[18])
         );
  DFFARX1 wdata_1_reg_17_ ( .D(N610), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[17])
         );
  DFFARX1 wdata_1_reg_16_ ( .D(N609), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[16])
         );
  DFFARX1 wdata_1_reg_15_ ( .D(N608), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[15])
         );
  DFFARX1 wdata_1_reg_14_ ( .D(N607), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[14])
         );
  DFFARX1 wdata_1_reg_13_ ( .D(N606), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[13])
         );
  DFFARX1 wdata_1_reg_12_ ( .D(N605), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[12])
         );
  DFFARX1 wdata_1_reg_11_ ( .D(N604), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[11])
         );
  DFFARX1 wdata_1_reg_10_ ( .D(N603), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[10])
         );
  DFFARX1 wdata_1_reg_9_ ( .D(N602), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[9])
         );
  DFFARX1 wdata_1_reg_8_ ( .D(N601), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[8])
         );
  DFFARX1 wdata_1_reg_7_ ( .D(N600), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[7])
         );
  DFFARX1 wdata_1_reg_6_ ( .D(N599), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[6])
         );
  DFFARX1 wdata_1_reg_5_ ( .D(N598), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[5])
         );
  DFFARX1 wdata_1_reg_4_ ( .D(N597), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[4])
         );
  DFFARX1 wdata_1_reg_3_ ( .D(N596), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[3])
         );
  DFFARX1 wdata_1_reg_2_ ( .D(N595), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[2])
         );
  DFFARX1 wdata_1_reg_1_ ( .D(N594), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[1])
         );
  DFFARX1 wdata_1_reg_0_ ( .D(N593), .CLK(clk), .RSTB(rst_n), .Q(wdata_1[0])
         );
  DFFARX1 wdata_0_reg_63_ ( .D(N720), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[63])
         );
  DFFARX1 wdata_0_reg_62_ ( .D(N719), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[62])
         );
  DFFARX1 wdata_0_reg_61_ ( .D(N718), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[61])
         );
  DFFARX1 wdata_0_reg_60_ ( .D(N717), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[60])
         );
  DFFARX1 wdata_0_reg_59_ ( .D(N716), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[59])
         );
  DFFARX1 wdata_0_reg_58_ ( .D(N715), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[58])
         );
  DFFARX1 wdata_0_reg_57_ ( .D(N714), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[57])
         );
  DFFARX1 wdata_0_reg_56_ ( .D(N713), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[56])
         );
  DFFARX1 wdata_0_reg_55_ ( .D(N712), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[55])
         );
  DFFARX1 wdata_0_reg_54_ ( .D(N711), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[54])
         );
  DFFARX1 wdata_0_reg_53_ ( .D(N710), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[53])
         );
  DFFARX1 wdata_0_reg_52_ ( .D(N709), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[52])
         );
  DFFARX1 wdata_0_reg_51_ ( .D(N708), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[51])
         );
  DFFARX1 wdata_0_reg_50_ ( .D(N707), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[50])
         );
  DFFARX1 wdata_0_reg_49_ ( .D(N706), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[49])
         );
  DFFARX1 wdata_0_reg_48_ ( .D(N705), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[48])
         );
  DFFARX1 wdata_0_reg_47_ ( .D(N704), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[47])
         );
  DFFARX1 wdata_0_reg_46_ ( .D(N703), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[46])
         );
  DFFARX1 wdata_0_reg_45_ ( .D(N702), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[45])
         );
  DFFARX1 wdata_0_reg_44_ ( .D(N701), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[44])
         );
  DFFARX1 wdata_0_reg_43_ ( .D(N700), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[43])
         );
  DFFARX1 wdata_0_reg_42_ ( .D(N699), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[42])
         );
  DFFARX1 wdata_0_reg_41_ ( .D(N698), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[41])
         );
  DFFARX1 wdata_0_reg_40_ ( .D(N697), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[40])
         );
  DFFARX1 wdata_0_reg_39_ ( .D(N696), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[39])
         );
  DFFARX1 wdata_0_reg_38_ ( .D(N695), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[38])
         );
  DFFARX1 wdata_0_reg_37_ ( .D(N694), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[37])
         );
  DFFARX1 wdata_0_reg_36_ ( .D(N693), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[36])
         );
  DFFARX1 wdata_0_reg_35_ ( .D(N692), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[35])
         );
  DFFARX1 wdata_0_reg_34_ ( .D(N691), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[34])
         );
  DFFARX1 wdata_0_reg_33_ ( .D(N690), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[33])
         );
  DFFARX1 wdata_0_reg_32_ ( .D(N689), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[32])
         );
  DFFARX1 wdata_0_reg_31_ ( .D(N688), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[31])
         );
  DFFARX1 wdata_0_reg_30_ ( .D(N687), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[30])
         );
  DFFARX1 wdata_0_reg_29_ ( .D(N686), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[29])
         );
  DFFARX1 wdata_0_reg_28_ ( .D(N685), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[28])
         );
  DFFARX1 wdata_0_reg_27_ ( .D(N684), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[27])
         );
  DFFARX1 wdata_0_reg_26_ ( .D(N683), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[26])
         );
  DFFARX1 wdata_0_reg_25_ ( .D(N682), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[25])
         );
  DFFARX1 wdata_0_reg_24_ ( .D(N681), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[24])
         );
  DFFARX1 wdata_0_reg_23_ ( .D(N680), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[23])
         );
  DFFARX1 wdata_0_reg_22_ ( .D(N679), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[22])
         );
  DFFARX1 wdata_0_reg_21_ ( .D(N678), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[21])
         );
  DFFARX1 wdata_0_reg_20_ ( .D(N677), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[20])
         );
  DFFARX1 wdata_0_reg_19_ ( .D(N676), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[19])
         );
  DFFARX1 wdata_0_reg_18_ ( .D(N675), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[18])
         );
  DFFARX1 wdata_0_reg_17_ ( .D(N674), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[17])
         );
  DFFARX1 wdata_0_reg_16_ ( .D(N673), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[16])
         );
  DFFARX1 wdata_0_reg_15_ ( .D(N672), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[15])
         );
  DFFARX1 wdata_0_reg_14_ ( .D(N671), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[14])
         );
  DFFARX1 wdata_0_reg_13_ ( .D(N670), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[13])
         );
  DFFARX1 wdata_0_reg_12_ ( .D(N669), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[12])
         );
  DFFARX1 wdata_0_reg_11_ ( .D(N668), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[11])
         );
  DFFARX1 wdata_0_reg_10_ ( .D(N667), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[10])
         );
  DFFARX1 wdata_0_reg_9_ ( .D(N666), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[9])
         );
  DFFARX1 wdata_0_reg_8_ ( .D(N665), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[8])
         );
  DFFARX1 wdata_0_reg_7_ ( .D(N664), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[7])
         );
  DFFARX1 wdata_0_reg_6_ ( .D(N663), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[6])
         );
  DFFARX1 wdata_0_reg_5_ ( .D(N662), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[5])
         );
  DFFARX1 wdata_0_reg_4_ ( .D(N661), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[4])
         );
  DFFARX1 wdata_0_reg_3_ ( .D(N660), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[3])
         );
  DFFARX1 wdata_0_reg_2_ ( .D(N659), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[2])
         );
  DFFARX1 wdata_0_reg_1_ ( .D(N658), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[1])
         );
  DFFARX1 wdata_0_reg_0_ ( .D(N657), .CLK(clk), .RSTB(rst_n), .Q(wdata_0[0])
         );
  DFFARX1 address_7_reg_15_ ( .D(N96), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[15]) );
  DFFARX1 address_7_reg_14_ ( .D(N95), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[14]) );
  DFFARX1 address_7_reg_13_ ( .D(N94), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[13]) );
  DFFARX1 address_7_reg_12_ ( .D(N93), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[12]) );
  DFFARX1 address_7_reg_11_ ( .D(N92), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[11]) );
  DFFARX1 address_7_reg_10_ ( .D(N91), .CLK(clk), .RSTB(rst_n), .Q(
        address_7[10]) );
  DFFARX1 address_7_reg_9_ ( .D(N90), .CLK(clk), .RSTB(rst_n), .Q(address_7[9]) );
  DFFARX1 address_7_reg_8_ ( .D(N89), .CLK(clk), .RSTB(rst_n), .Q(address_7[8]) );
  DFFARX1 address_7_reg_7_ ( .D(N88), .CLK(clk), .RSTB(rst_n), .Q(address_7[7]) );
  DFFARX1 address_7_reg_6_ ( .D(N87), .CLK(clk), .RSTB(rst_n), .Q(address_7[6]) );
  DFFARX1 address_7_reg_5_ ( .D(N86), .CLK(clk), .RSTB(rst_n), .Q(address_7[5]) );
  DFFARX1 address_7_reg_4_ ( .D(N85), .CLK(clk), .RSTB(rst_n), .Q(address_7[4]) );
  DFFARX1 address_7_reg_3_ ( .D(N84), .CLK(clk), .RSTB(rst_n), .Q(address_7[3]) );
  DFFARX1 address_7_reg_2_ ( .D(N83), .CLK(clk), .RSTB(rst_n), .Q(address_7[2]) );
  DFFARX1 address_7_reg_1_ ( .D(N82), .CLK(clk), .RSTB(rst_n), .Q(address_7[1]) );
  DFFARX1 address_7_reg_0_ ( .D(N81), .CLK(clk), .RSTB(rst_n), .Q(address_7[0]) );
  DFFARX1 address_6_reg_15_ ( .D(N112), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[15]) );
  DFFARX1 address_6_reg_14_ ( .D(N111), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[14]) );
  DFFARX1 address_6_reg_13_ ( .D(N110), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[13]) );
  DFFARX1 address_6_reg_12_ ( .D(N109), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[12]) );
  DFFARX1 address_6_reg_11_ ( .D(N108), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[11]) );
  DFFARX1 address_6_reg_10_ ( .D(N107), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[10]) );
  DFFARX1 address_6_reg_9_ ( .D(N106), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[9]) );
  DFFARX1 address_6_reg_8_ ( .D(N105), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[8]) );
  DFFARX1 address_6_reg_7_ ( .D(N104), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[7]) );
  DFFARX1 address_6_reg_6_ ( .D(N103), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[6]) );
  DFFARX1 address_6_reg_5_ ( .D(N102), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[5]) );
  DFFARX1 address_6_reg_4_ ( .D(N101), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[4]) );
  DFFARX1 address_6_reg_3_ ( .D(N100), .CLK(clk), .RSTB(rst_n), .Q(
        address_6[3]) );
  DFFARX1 address_6_reg_2_ ( .D(N99), .CLK(clk), .RSTB(rst_n), .Q(address_6[2]) );
  DFFARX1 address_6_reg_1_ ( .D(N98), .CLK(clk), .RSTB(rst_n), .Q(address_6[1]) );
  DFFARX1 address_6_reg_0_ ( .D(N97), .CLK(clk), .RSTB(rst_n), .Q(address_6[0]) );
  DFFARX1 address_5_reg_15_ ( .D(N128), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[15]) );
  DFFARX1 address_5_reg_14_ ( .D(N127), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[14]) );
  DFFARX1 address_5_reg_13_ ( .D(N126), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[13]) );
  DFFARX1 address_5_reg_12_ ( .D(N125), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[12]) );
  DFFARX1 address_5_reg_11_ ( .D(N124), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[11]) );
  DFFARX1 address_5_reg_10_ ( .D(N123), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[10]) );
  DFFARX1 address_5_reg_9_ ( .D(N122), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[9]) );
  DFFARX1 address_5_reg_8_ ( .D(N121), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[8]) );
  DFFARX1 address_5_reg_7_ ( .D(N120), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[7]) );
  DFFARX1 address_5_reg_6_ ( .D(N119), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[6]) );
  DFFARX1 address_5_reg_5_ ( .D(N118), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[5]) );
  DFFARX1 address_5_reg_4_ ( .D(N117), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[4]) );
  DFFARX1 address_5_reg_3_ ( .D(N116), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[3]) );
  DFFARX1 address_5_reg_2_ ( .D(N115), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[2]) );
  DFFARX1 address_5_reg_1_ ( .D(N114), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[1]) );
  DFFARX1 address_5_reg_0_ ( .D(N113), .CLK(clk), .RSTB(rst_n), .Q(
        address_5[0]) );
  NOR2X0 U93 ( .IN1(n713), .IN2(n800), .QN(N99) );
  NOR2X0 U94 ( .IN1(n713), .IN2(n801), .QN(N98) );
  NOR2X0 U95 ( .IN1(n713), .IN2(n802), .QN(N97) );
  NOR2X0 U96 ( .IN1(n803), .IN2(n787), .QN(N96) );
  NOR2X0 U97 ( .IN1(n803), .IN2(n788), .QN(N95) );
  NOR2X0 U98 ( .IN1(n803), .IN2(n789), .QN(N94) );
  NOR2X0 U99 ( .IN1(n803), .IN2(n790), .QN(N93) );
  NOR2X0 U100 ( .IN1(n803), .IN2(n791), .QN(N92) );
  NOR2X0 U101 ( .IN1(n803), .IN2(n792), .QN(N91) );
  NOR2X0 U102 ( .IN1(n803), .IN2(n793), .QN(N90) );
  NOR2X0 U103 ( .IN1(n803), .IN2(n794), .QN(N89) );
  NOR2X0 U104 ( .IN1(n803), .IN2(n795), .QN(N88) );
  NOR2X0 U105 ( .IN1(n803), .IN2(n796), .QN(N87) );
  NOR2X0 U106 ( .IN1(n803), .IN2(n797), .QN(N86) );
  NOR2X0 U107 ( .IN1(n803), .IN2(n798), .QN(N85) );
  NOR2X0 U108 ( .IN1(n803), .IN2(n799), .QN(N84) );
  NOR2X0 U109 ( .IN1(n803), .IN2(n800), .QN(N83) );
  NOR2X0 U110 ( .IN1(n803), .IN2(n801), .QN(N82) );
  NOR2X0 U111 ( .IN1(n803), .IN2(n802), .QN(N81) );
  OR2X1 U112 ( .IN1(n804), .IN2(n805), .Q(N79) );
  AO221X1 U113 ( .IN1(n806), .IN2(rdata_1[63]), .IN3(n807), .IN4(rdata_0[63]), 
        .IN5(n808), .Q(n805) );
  AO22X1 U114 ( .IN1(n809), .IN2(rdata_2[63]), .IN3(n720), .IN4(rdata_7[63]), 
        .Q(n808) );
  AO221X1 U115 ( .IN1(n810), .IN2(rdata_4[63]), .IN3(n811), .IN4(rdata_3[63]), 
        .IN5(n812), .Q(n804) );
  AO22X1 U116 ( .IN1(n813), .IN2(rdata_5[63]), .IN3(n814), .IN4(rdata_6[63]), 
        .Q(n812) );
  OR2X1 U117 ( .IN1(n815), .IN2(n816), .Q(N78) );
  AO221X1 U118 ( .IN1(n806), .IN2(rdata_1[62]), .IN3(n807), .IN4(rdata_0[62]), 
        .IN5(n817), .Q(n816) );
  AO22X1 U119 ( .IN1(n809), .IN2(rdata_2[62]), .IN3(n720), .IN4(rdata_7[62]), 
        .Q(n817) );
  AO221X1 U120 ( .IN1(n810), .IN2(rdata_4[62]), .IN3(n811), .IN4(rdata_3[62]), 
        .IN5(n818), .Q(n815) );
  AO22X1 U121 ( .IN1(n813), .IN2(rdata_5[62]), .IN3(n814), .IN4(rdata_6[62]), 
        .Q(n818) );
  OR2X1 U122 ( .IN1(n819), .IN2(n820), .Q(N77) );
  AO221X1 U123 ( .IN1(n806), .IN2(rdata_1[61]), .IN3(n807), .IN4(rdata_0[61]), 
        .IN5(n821), .Q(n820) );
  AO22X1 U124 ( .IN1(n809), .IN2(rdata_2[61]), .IN3(n720), .IN4(rdata_7[61]), 
        .Q(n821) );
  AO221X1 U125 ( .IN1(n810), .IN2(rdata_4[61]), .IN3(n811), .IN4(rdata_3[61]), 
        .IN5(n822), .Q(n819) );
  AO22X1 U126 ( .IN1(n813), .IN2(rdata_5[61]), .IN3(n814), .IN4(rdata_6[61]), 
        .Q(n822) );
  OR2X1 U127 ( .IN1(n823), .IN2(n824), .Q(N76) );
  AO221X1 U128 ( .IN1(n806), .IN2(rdata_1[60]), .IN3(n807), .IN4(rdata_0[60]), 
        .IN5(n825), .Q(n824) );
  AO22X1 U129 ( .IN1(n809), .IN2(rdata_2[60]), .IN3(n720), .IN4(rdata_7[60]), 
        .Q(n825) );
  AO221X1 U130 ( .IN1(n810), .IN2(rdata_4[60]), .IN3(n811), .IN4(rdata_3[60]), 
        .IN5(n826), .Q(n823) );
  AO22X1 U131 ( .IN1(n813), .IN2(rdata_5[60]), .IN3(n814), .IN4(rdata_6[60]), 
        .Q(n826) );
  OR2X1 U132 ( .IN1(n827), .IN2(n828), .Q(N75) );
  AO221X1 U133 ( .IN1(n806), .IN2(rdata_1[59]), .IN3(n807), .IN4(rdata_0[59]), 
        .IN5(n829), .Q(n828) );
  AO22X1 U134 ( .IN1(n809), .IN2(rdata_2[59]), .IN3(n720), .IN4(rdata_7[59]), 
        .Q(n829) );
  AO221X1 U135 ( .IN1(n810), .IN2(rdata_4[59]), .IN3(n811), .IN4(rdata_3[59]), 
        .IN5(n830), .Q(n827) );
  AO22X1 U136 ( .IN1(n813), .IN2(rdata_5[59]), .IN3(n814), .IN4(rdata_6[59]), 
        .Q(n830) );
  OR2X1 U137 ( .IN1(n831), .IN2(n832), .Q(N74) );
  AO221X1 U138 ( .IN1(n806), .IN2(rdata_1[58]), .IN3(n807), .IN4(rdata_0[58]), 
        .IN5(n833), .Q(n832) );
  AO22X1 U139 ( .IN1(n809), .IN2(rdata_2[58]), .IN3(n720), .IN4(rdata_7[58]), 
        .Q(n833) );
  AO221X1 U140 ( .IN1(n810), .IN2(rdata_4[58]), .IN3(n811), .IN4(rdata_3[58]), 
        .IN5(n834), .Q(n831) );
  AO22X1 U141 ( .IN1(n813), .IN2(rdata_5[58]), .IN3(n814), .IN4(rdata_6[58]), 
        .Q(n834) );
  OR2X1 U142 ( .IN1(n835), .IN2(n836), .Q(N73) );
  AO221X1 U143 ( .IN1(n806), .IN2(rdata_1[57]), .IN3(n807), .IN4(rdata_0[57]), 
        .IN5(n837), .Q(n836) );
  AO22X1 U144 ( .IN1(n809), .IN2(rdata_2[57]), .IN3(n720), .IN4(rdata_7[57]), 
        .Q(n837) );
  AO221X1 U145 ( .IN1(n810), .IN2(rdata_4[57]), .IN3(n811), .IN4(rdata_3[57]), 
        .IN5(n838), .Q(n835) );
  AO22X1 U146 ( .IN1(n813), .IN2(rdata_5[57]), .IN3(n814), .IN4(rdata_6[57]), 
        .Q(n838) );
  NOR2X0 U147 ( .IN1(n718), .IN2(n722), .QN(N728) );
  NOR2X0 U148 ( .IN1(n719), .IN2(n722), .QN(N727) );
  NOR2X0 U149 ( .IN1(n717), .IN2(n722), .QN(N726) );
  NOR2X0 U150 ( .IN1(n715), .IN2(n722), .QN(N725) );
  NOR2X0 U151 ( .IN1(n716), .IN2(n722), .QN(N724) );
  NOR2X0 U152 ( .IN1(n714), .IN2(n722), .QN(N723) );
  NOR2X0 U153 ( .IN1(n713), .IN2(n722), .QN(N722) );
  NOR2X0 U154 ( .IN1(n803), .IN2(n722), .QN(N721) );
  NOR2X0 U155 ( .IN1(n718), .IN2(n723), .QN(N720) );
  OR2X1 U156 ( .IN1(n839), .IN2(n840), .Q(N72) );
  AO221X1 U157 ( .IN1(n806), .IN2(rdata_1[56]), .IN3(n807), .IN4(rdata_0[56]), 
        .IN5(n841), .Q(n840) );
  AO22X1 U158 ( .IN1(n809), .IN2(rdata_2[56]), .IN3(n720), .IN4(rdata_7[56]), 
        .Q(n841) );
  AO221X1 U159 ( .IN1(n810), .IN2(rdata_4[56]), .IN3(n811), .IN4(rdata_3[56]), 
        .IN5(n842), .Q(n839) );
  AO22X1 U160 ( .IN1(n813), .IN2(rdata_5[56]), .IN3(n814), .IN4(rdata_6[56]), 
        .Q(n842) );
  NOR2X0 U161 ( .IN1(n718), .IN2(n724), .QN(N719) );
  NOR2X0 U162 ( .IN1(n718), .IN2(n725), .QN(N718) );
  NOR2X0 U163 ( .IN1(n718), .IN2(n726), .QN(N717) );
  NOR2X0 U164 ( .IN1(n718), .IN2(n727), .QN(N716) );
  NOR2X0 U165 ( .IN1(n718), .IN2(n728), .QN(N715) );
  NOR2X0 U166 ( .IN1(n718), .IN2(n729), .QN(N714) );
  NOR2X0 U167 ( .IN1(n718), .IN2(n730), .QN(N713) );
  NOR2X0 U168 ( .IN1(n718), .IN2(n731), .QN(N712) );
  NOR2X0 U169 ( .IN1(n718), .IN2(n732), .QN(N711) );
  NOR2X0 U170 ( .IN1(n718), .IN2(n733), .QN(N710) );
  OR2X1 U171 ( .IN1(n843), .IN2(n844), .Q(N71) );
  AO221X1 U172 ( .IN1(n806), .IN2(rdata_1[55]), .IN3(n807), .IN4(rdata_0[55]), 
        .IN5(n845), .Q(n844) );
  AO22X1 U173 ( .IN1(n809), .IN2(rdata_2[55]), .IN3(n720), .IN4(rdata_7[55]), 
        .Q(n845) );
  AO221X1 U174 ( .IN1(n810), .IN2(rdata_4[55]), .IN3(n811), .IN4(rdata_3[55]), 
        .IN5(n846), .Q(n843) );
  AO22X1 U175 ( .IN1(n813), .IN2(rdata_5[55]), .IN3(n814), .IN4(rdata_6[55]), 
        .Q(n846) );
  NOR2X0 U176 ( .IN1(n718), .IN2(n734), .QN(N709) );
  NOR2X0 U177 ( .IN1(n718), .IN2(n735), .QN(N708) );
  NOR2X0 U178 ( .IN1(n718), .IN2(n736), .QN(N707) );
  NOR2X0 U179 ( .IN1(n718), .IN2(n737), .QN(N706) );
  NOR2X0 U180 ( .IN1(n718), .IN2(n738), .QN(N705) );
  NOR2X0 U181 ( .IN1(n718), .IN2(n739), .QN(N704) );
  NOR2X0 U182 ( .IN1(n718), .IN2(n740), .QN(N703) );
  NOR2X0 U183 ( .IN1(n718), .IN2(n741), .QN(N702) );
  NOR2X0 U184 ( .IN1(n718), .IN2(n742), .QN(N701) );
  NOR2X0 U185 ( .IN1(n718), .IN2(n743), .QN(N700) );
  OR2X1 U186 ( .IN1(n847), .IN2(n848), .Q(N70) );
  AO221X1 U187 ( .IN1(n806), .IN2(rdata_1[54]), .IN3(n807), .IN4(rdata_0[54]), 
        .IN5(n849), .Q(n848) );
  AO22X1 U188 ( .IN1(n809), .IN2(rdata_2[54]), .IN3(n720), .IN4(rdata_7[54]), 
        .Q(n849) );
  AO221X1 U189 ( .IN1(n810), .IN2(rdata_4[54]), .IN3(n811), .IN4(rdata_3[54]), 
        .IN5(n850), .Q(n847) );
  AO22X1 U190 ( .IN1(n813), .IN2(rdata_5[54]), .IN3(n814), .IN4(rdata_6[54]), 
        .Q(n850) );
  NOR2X0 U191 ( .IN1(n718), .IN2(n744), .QN(N699) );
  NOR2X0 U192 ( .IN1(n718), .IN2(n745), .QN(N698) );
  NOR2X0 U193 ( .IN1(n718), .IN2(n746), .QN(N697) );
  NOR2X0 U194 ( .IN1(n718), .IN2(n747), .QN(N696) );
  NOR2X0 U195 ( .IN1(n718), .IN2(n748), .QN(N695) );
  NOR2X0 U196 ( .IN1(n718), .IN2(n749), .QN(N694) );
  NOR2X0 U197 ( .IN1(n718), .IN2(n750), .QN(N693) );
  NOR2X0 U198 ( .IN1(n718), .IN2(n751), .QN(N692) );
  NOR2X0 U199 ( .IN1(n718), .IN2(n752), .QN(N691) );
  NOR2X0 U200 ( .IN1(n718), .IN2(n753), .QN(N690) );
  OR2X1 U201 ( .IN1(n851), .IN2(n852), .Q(N69) );
  AO221X1 U202 ( .IN1(n806), .IN2(rdata_1[53]), .IN3(n807), .IN4(rdata_0[53]), 
        .IN5(n853), .Q(n852) );
  AO22X1 U203 ( .IN1(n809), .IN2(rdata_2[53]), .IN3(n720), .IN4(rdata_7[53]), 
        .Q(n853) );
  AO221X1 U204 ( .IN1(n810), .IN2(rdata_4[53]), .IN3(n811), .IN4(rdata_3[53]), 
        .IN5(n854), .Q(n851) );
  AO22X1 U205 ( .IN1(n813), .IN2(rdata_5[53]), .IN3(n814), .IN4(rdata_6[53]), 
        .Q(n854) );
  NOR2X0 U206 ( .IN1(n718), .IN2(n754), .QN(N689) );
  NOR2X0 U207 ( .IN1(n718), .IN2(n755), .QN(N688) );
  NOR2X0 U208 ( .IN1(n718), .IN2(n756), .QN(N687) );
  NOR2X0 U209 ( .IN1(n718), .IN2(n757), .QN(N686) );
  NOR2X0 U210 ( .IN1(n718), .IN2(n758), .QN(N685) );
  NOR2X0 U211 ( .IN1(n718), .IN2(n759), .QN(N684) );
  NOR2X0 U212 ( .IN1(n718), .IN2(n760), .QN(N683) );
  NOR2X0 U213 ( .IN1(n718), .IN2(n761), .QN(N682) );
  NOR2X0 U214 ( .IN1(n718), .IN2(n762), .QN(N681) );
  NOR2X0 U215 ( .IN1(n718), .IN2(n763), .QN(N680) );
  OR2X1 U216 ( .IN1(n855), .IN2(n856), .Q(N68) );
  AO221X1 U217 ( .IN1(n806), .IN2(rdata_1[52]), .IN3(n807), .IN4(rdata_0[52]), 
        .IN5(n857), .Q(n856) );
  AO22X1 U218 ( .IN1(n809), .IN2(rdata_2[52]), .IN3(n720), .IN4(rdata_7[52]), 
        .Q(n857) );
  AO221X1 U219 ( .IN1(n810), .IN2(rdata_4[52]), .IN3(n811), .IN4(rdata_3[52]), 
        .IN5(n858), .Q(n855) );
  AO22X1 U220 ( .IN1(n813), .IN2(rdata_5[52]), .IN3(n814), .IN4(rdata_6[52]), 
        .Q(n858) );
  NOR2X0 U221 ( .IN1(n718), .IN2(n764), .QN(N679) );
  NOR2X0 U222 ( .IN1(n718), .IN2(n765), .QN(N678) );
  NOR2X0 U223 ( .IN1(n718), .IN2(n766), .QN(N677) );
  NOR2X0 U224 ( .IN1(n718), .IN2(n767), .QN(N676) );
  NOR2X0 U225 ( .IN1(n718), .IN2(n768), .QN(N675) );
  NOR2X0 U226 ( .IN1(n718), .IN2(n769), .QN(N674) );
  NOR2X0 U227 ( .IN1(n718), .IN2(n770), .QN(N673) );
  NOR2X0 U228 ( .IN1(n718), .IN2(n771), .QN(N672) );
  NOR2X0 U229 ( .IN1(n718), .IN2(n772), .QN(N671) );
  NOR2X0 U230 ( .IN1(n718), .IN2(n773), .QN(N670) );
  OR2X1 U231 ( .IN1(n859), .IN2(n860), .Q(N67) );
  AO221X1 U232 ( .IN1(n806), .IN2(rdata_1[51]), .IN3(n807), .IN4(rdata_0[51]), 
        .IN5(n861), .Q(n860) );
  AO22X1 U233 ( .IN1(n809), .IN2(rdata_2[51]), .IN3(n720), .IN4(rdata_7[51]), 
        .Q(n861) );
  AO221X1 U234 ( .IN1(n810), .IN2(rdata_4[51]), .IN3(n811), .IN4(rdata_3[51]), 
        .IN5(n862), .Q(n859) );
  AO22X1 U235 ( .IN1(n813), .IN2(rdata_5[51]), .IN3(n814), .IN4(rdata_6[51]), 
        .Q(n862) );
  NOR2X0 U236 ( .IN1(n718), .IN2(n774), .QN(N669) );
  NOR2X0 U237 ( .IN1(n718), .IN2(n775), .QN(N668) );
  NOR2X0 U238 ( .IN1(n718), .IN2(n776), .QN(N667) );
  NOR2X0 U239 ( .IN1(n718), .IN2(n777), .QN(N666) );
  NOR2X0 U240 ( .IN1(n718), .IN2(n778), .QN(N665) );
  NOR2X0 U241 ( .IN1(n718), .IN2(n779), .QN(N664) );
  NOR2X0 U242 ( .IN1(n718), .IN2(n780), .QN(N663) );
  NOR2X0 U243 ( .IN1(n718), .IN2(n781), .QN(N662) );
  NOR2X0 U244 ( .IN1(n718), .IN2(n782), .QN(N661) );
  NOR2X0 U245 ( .IN1(n718), .IN2(n783), .QN(N660) );
  OR2X1 U246 ( .IN1(n863), .IN2(n864), .Q(N66) );
  AO221X1 U247 ( .IN1(n806), .IN2(rdata_1[50]), .IN3(n807), .IN4(rdata_0[50]), 
        .IN5(n865), .Q(n864) );
  AO22X1 U248 ( .IN1(n809), .IN2(rdata_2[50]), .IN3(n720), .IN4(rdata_7[50]), 
        .Q(n865) );
  AO221X1 U249 ( .IN1(n810), .IN2(rdata_4[50]), .IN3(n811), .IN4(rdata_3[50]), 
        .IN5(n866), .Q(n863) );
  AO22X1 U250 ( .IN1(n813), .IN2(rdata_5[50]), .IN3(n814), .IN4(rdata_6[50]), 
        .Q(n866) );
  NOR2X0 U251 ( .IN1(n718), .IN2(n784), .QN(N659) );
  NOR2X0 U252 ( .IN1(n718), .IN2(n785), .QN(N658) );
  NOR2X0 U253 ( .IN1(n718), .IN2(n786), .QN(N657) );
  NOR2X0 U254 ( .IN1(n719), .IN2(n723), .QN(N656) );
  NOR2X0 U255 ( .IN1(n719), .IN2(n724), .QN(N655) );
  NOR2X0 U256 ( .IN1(n719), .IN2(n725), .QN(N654) );
  NOR2X0 U257 ( .IN1(n719), .IN2(n726), .QN(N653) );
  NOR2X0 U258 ( .IN1(n719), .IN2(n727), .QN(N652) );
  NOR2X0 U259 ( .IN1(n719), .IN2(n728), .QN(N651) );
  NOR2X0 U260 ( .IN1(n719), .IN2(n729), .QN(N650) );
  OR2X1 U261 ( .IN1(n867), .IN2(n868), .Q(N65) );
  AO221X1 U262 ( .IN1(n806), .IN2(rdata_1[49]), .IN3(n807), .IN4(rdata_0[49]), 
        .IN5(n869), .Q(n868) );
  AO22X1 U263 ( .IN1(n809), .IN2(rdata_2[49]), .IN3(n720), .IN4(rdata_7[49]), 
        .Q(n869) );
  AO221X1 U264 ( .IN1(n810), .IN2(rdata_4[49]), .IN3(n811), .IN4(rdata_3[49]), 
        .IN5(n870), .Q(n867) );
  AO22X1 U265 ( .IN1(n813), .IN2(rdata_5[49]), .IN3(n814), .IN4(rdata_6[49]), 
        .Q(n870) );
  NOR2X0 U266 ( .IN1(n719), .IN2(n730), .QN(N649) );
  NOR2X0 U267 ( .IN1(n719), .IN2(n731), .QN(N648) );
  NOR2X0 U268 ( .IN1(n719), .IN2(n732), .QN(N647) );
  NOR2X0 U269 ( .IN1(n719), .IN2(n733), .QN(N646) );
  NOR2X0 U270 ( .IN1(n719), .IN2(n734), .QN(N645) );
  NOR2X0 U271 ( .IN1(n719), .IN2(n735), .QN(N644) );
  NOR2X0 U272 ( .IN1(n719), .IN2(n736), .QN(N643) );
  NOR2X0 U273 ( .IN1(n719), .IN2(n737), .QN(N642) );
  NOR2X0 U274 ( .IN1(n719), .IN2(n738), .QN(N641) );
  NOR2X0 U275 ( .IN1(n719), .IN2(n739), .QN(N640) );
  OR2X1 U276 ( .IN1(n871), .IN2(n872), .Q(N64) );
  AO221X1 U277 ( .IN1(n806), .IN2(rdata_1[48]), .IN3(n807), .IN4(rdata_0[48]), 
        .IN5(n873), .Q(n872) );
  AO22X1 U278 ( .IN1(n809), .IN2(rdata_2[48]), .IN3(n720), .IN4(rdata_7[48]), 
        .Q(n873) );
  AO221X1 U279 ( .IN1(n810), .IN2(rdata_4[48]), .IN3(n811), .IN4(rdata_3[48]), 
        .IN5(n874), .Q(n871) );
  AO22X1 U280 ( .IN1(n813), .IN2(rdata_5[48]), .IN3(n814), .IN4(rdata_6[48]), 
        .Q(n874) );
  NOR2X0 U281 ( .IN1(n719), .IN2(n740), .QN(N639) );
  NOR2X0 U282 ( .IN1(n719), .IN2(n741), .QN(N638) );
  NOR2X0 U283 ( .IN1(n719), .IN2(n742), .QN(N637) );
  NOR2X0 U284 ( .IN1(n719), .IN2(n743), .QN(N636) );
  NOR2X0 U285 ( .IN1(n719), .IN2(n744), .QN(N635) );
  NOR2X0 U286 ( .IN1(n719), .IN2(n745), .QN(N634) );
  NOR2X0 U287 ( .IN1(n719), .IN2(n746), .QN(N633) );
  NOR2X0 U288 ( .IN1(n719), .IN2(n747), .QN(N632) );
  NOR2X0 U289 ( .IN1(n719), .IN2(n748), .QN(N631) );
  NOR2X0 U290 ( .IN1(n719), .IN2(n749), .QN(N630) );
  OR2X1 U291 ( .IN1(n875), .IN2(n876), .Q(N63) );
  AO221X1 U292 ( .IN1(n806), .IN2(rdata_1[47]), .IN3(n807), .IN4(rdata_0[47]), 
        .IN5(n877), .Q(n876) );
  AO22X1 U293 ( .IN1(n809), .IN2(rdata_2[47]), .IN3(n720), .IN4(rdata_7[47]), 
        .Q(n877) );
  AO221X1 U294 ( .IN1(n810), .IN2(rdata_4[47]), .IN3(n811), .IN4(rdata_3[47]), 
        .IN5(n878), .Q(n875) );
  AO22X1 U295 ( .IN1(n813), .IN2(rdata_5[47]), .IN3(n814), .IN4(rdata_6[47]), 
        .Q(n878) );
  NOR2X0 U296 ( .IN1(n719), .IN2(n750), .QN(N629) );
  NOR2X0 U297 ( .IN1(n719), .IN2(n751), .QN(N628) );
  NOR2X0 U298 ( .IN1(n719), .IN2(n752), .QN(N627) );
  NOR2X0 U299 ( .IN1(n719), .IN2(n753), .QN(N626) );
  NOR2X0 U300 ( .IN1(n719), .IN2(n754), .QN(N625) );
  NOR2X0 U301 ( .IN1(n719), .IN2(n755), .QN(N624) );
  NOR2X0 U302 ( .IN1(n719), .IN2(n756), .QN(N623) );
  NOR2X0 U303 ( .IN1(n719), .IN2(n757), .QN(N622) );
  NOR2X0 U304 ( .IN1(n719), .IN2(n758), .QN(N621) );
  NOR2X0 U305 ( .IN1(n719), .IN2(n759), .QN(N620) );
  OR2X1 U306 ( .IN1(n879), .IN2(n880), .Q(N62) );
  AO221X1 U307 ( .IN1(n806), .IN2(rdata_1[46]), .IN3(n807), .IN4(rdata_0[46]), 
        .IN5(n881), .Q(n880) );
  AO22X1 U308 ( .IN1(n809), .IN2(rdata_2[46]), .IN3(n720), .IN4(rdata_7[46]), 
        .Q(n881) );
  AO221X1 U309 ( .IN1(n810), .IN2(rdata_4[46]), .IN3(n811), .IN4(rdata_3[46]), 
        .IN5(n882), .Q(n879) );
  AO22X1 U310 ( .IN1(n813), .IN2(rdata_5[46]), .IN3(n814), .IN4(rdata_6[46]), 
        .Q(n882) );
  NOR2X0 U311 ( .IN1(n719), .IN2(n760), .QN(N619) );
  NOR2X0 U312 ( .IN1(n719), .IN2(n761), .QN(N618) );
  NOR2X0 U313 ( .IN1(n719), .IN2(n762), .QN(N617) );
  NOR2X0 U314 ( .IN1(n719), .IN2(n763), .QN(N616) );
  NOR2X0 U315 ( .IN1(n719), .IN2(n764), .QN(N615) );
  NOR2X0 U316 ( .IN1(n719), .IN2(n765), .QN(N614) );
  NOR2X0 U317 ( .IN1(n719), .IN2(n766), .QN(N613) );
  NOR2X0 U318 ( .IN1(n719), .IN2(n767), .QN(N612) );
  NOR2X0 U319 ( .IN1(n719), .IN2(n768), .QN(N611) );
  NOR2X0 U320 ( .IN1(n719), .IN2(n769), .QN(N610) );
  OR2X1 U321 ( .IN1(n883), .IN2(n884), .Q(N61) );
  AO221X1 U322 ( .IN1(n806), .IN2(rdata_1[45]), .IN3(n807), .IN4(rdata_0[45]), 
        .IN5(n885), .Q(n884) );
  AO22X1 U323 ( .IN1(n809), .IN2(rdata_2[45]), .IN3(n720), .IN4(rdata_7[45]), 
        .Q(n885) );
  AO221X1 U324 ( .IN1(n810), .IN2(rdata_4[45]), .IN3(n811), .IN4(rdata_3[45]), 
        .IN5(n886), .Q(n883) );
  AO22X1 U325 ( .IN1(n813), .IN2(rdata_5[45]), .IN3(n814), .IN4(rdata_6[45]), 
        .Q(n886) );
  NOR2X0 U326 ( .IN1(n719), .IN2(n770), .QN(N609) );
  NOR2X0 U327 ( .IN1(n719), .IN2(n771), .QN(N608) );
  NOR2X0 U328 ( .IN1(n719), .IN2(n772), .QN(N607) );
  NOR2X0 U329 ( .IN1(n719), .IN2(n773), .QN(N606) );
  NOR2X0 U330 ( .IN1(n719), .IN2(n774), .QN(N605) );
  NOR2X0 U331 ( .IN1(n719), .IN2(n775), .QN(N604) );
  NOR2X0 U332 ( .IN1(n719), .IN2(n776), .QN(N603) );
  NOR2X0 U333 ( .IN1(n719), .IN2(n777), .QN(N602) );
  NOR2X0 U334 ( .IN1(n719), .IN2(n778), .QN(N601) );
  NOR2X0 U335 ( .IN1(n719), .IN2(n779), .QN(N600) );
  OR2X1 U336 ( .IN1(n887), .IN2(n888), .Q(N60) );
  AO221X1 U337 ( .IN1(n806), .IN2(rdata_1[44]), .IN3(n807), .IN4(rdata_0[44]), 
        .IN5(n889), .Q(n888) );
  AO22X1 U338 ( .IN1(n809), .IN2(rdata_2[44]), .IN3(n720), .IN4(rdata_7[44]), 
        .Q(n889) );
  AO221X1 U339 ( .IN1(n810), .IN2(rdata_4[44]), .IN3(n811), .IN4(rdata_3[44]), 
        .IN5(n890), .Q(n887) );
  AO22X1 U340 ( .IN1(n813), .IN2(rdata_5[44]), .IN3(n814), .IN4(rdata_6[44]), 
        .Q(n890) );
  NOR2X0 U341 ( .IN1(n719), .IN2(n780), .QN(N599) );
  NOR2X0 U342 ( .IN1(n719), .IN2(n781), .QN(N598) );
  NOR2X0 U343 ( .IN1(n719), .IN2(n782), .QN(N597) );
  NOR2X0 U344 ( .IN1(n719), .IN2(n783), .QN(N596) );
  NOR2X0 U345 ( .IN1(n719), .IN2(n784), .QN(N595) );
  NOR2X0 U346 ( .IN1(n719), .IN2(n785), .QN(N594) );
  NOR2X0 U347 ( .IN1(n719), .IN2(n786), .QN(N593) );
  NOR2X0 U348 ( .IN1(n717), .IN2(n723), .QN(N592) );
  NOR2X0 U349 ( .IN1(n717), .IN2(n724), .QN(N591) );
  NOR2X0 U350 ( .IN1(n717), .IN2(n725), .QN(N590) );
  OR2X1 U351 ( .IN1(n891), .IN2(n892), .Q(N59) );
  AO221X1 U352 ( .IN1(n806), .IN2(rdata_1[43]), .IN3(n807), .IN4(rdata_0[43]), 
        .IN5(n893), .Q(n892) );
  AO22X1 U353 ( .IN1(n809), .IN2(rdata_2[43]), .IN3(n720), .IN4(rdata_7[43]), 
        .Q(n893) );
  AO221X1 U354 ( .IN1(n810), .IN2(rdata_4[43]), .IN3(n811), .IN4(rdata_3[43]), 
        .IN5(n894), .Q(n891) );
  AO22X1 U355 ( .IN1(n813), .IN2(rdata_5[43]), .IN3(n814), .IN4(rdata_6[43]), 
        .Q(n894) );
  NOR2X0 U356 ( .IN1(n717), .IN2(n726), .QN(N589) );
  NOR2X0 U357 ( .IN1(n717), .IN2(n727), .QN(N588) );
  NOR2X0 U358 ( .IN1(n717), .IN2(n728), .QN(N587) );
  NOR2X0 U359 ( .IN1(n717), .IN2(n729), .QN(N586) );
  NOR2X0 U360 ( .IN1(n717), .IN2(n730), .QN(N585) );
  NOR2X0 U361 ( .IN1(n717), .IN2(n731), .QN(N584) );
  NOR2X0 U362 ( .IN1(n717), .IN2(n732), .QN(N583) );
  NOR2X0 U363 ( .IN1(n717), .IN2(n733), .QN(N582) );
  NOR2X0 U364 ( .IN1(n717), .IN2(n734), .QN(N581) );
  NOR2X0 U365 ( .IN1(n717), .IN2(n735), .QN(N580) );
  OR2X1 U366 ( .IN1(n895), .IN2(n896), .Q(N58) );
  AO221X1 U367 ( .IN1(n806), .IN2(rdata_1[42]), .IN3(n807), .IN4(rdata_0[42]), 
        .IN5(n897), .Q(n896) );
  AO22X1 U368 ( .IN1(n809), .IN2(rdata_2[42]), .IN3(n720), .IN4(rdata_7[42]), 
        .Q(n897) );
  AO221X1 U369 ( .IN1(n810), .IN2(rdata_4[42]), .IN3(n811), .IN4(rdata_3[42]), 
        .IN5(n898), .Q(n895) );
  AO22X1 U370 ( .IN1(n813), .IN2(rdata_5[42]), .IN3(n814), .IN4(rdata_6[42]), 
        .Q(n898) );
  NOR2X0 U371 ( .IN1(n717), .IN2(n736), .QN(N579) );
  NOR2X0 U372 ( .IN1(n717), .IN2(n737), .QN(N578) );
  NOR2X0 U373 ( .IN1(n717), .IN2(n738), .QN(N577) );
  NOR2X0 U374 ( .IN1(n717), .IN2(n739), .QN(N576) );
  NOR2X0 U375 ( .IN1(n717), .IN2(n740), .QN(N575) );
  NOR2X0 U376 ( .IN1(n717), .IN2(n741), .QN(N574) );
  NOR2X0 U377 ( .IN1(n717), .IN2(n742), .QN(N573) );
  NOR2X0 U378 ( .IN1(n717), .IN2(n743), .QN(N572) );
  NOR2X0 U379 ( .IN1(n717), .IN2(n744), .QN(N571) );
  NOR2X0 U380 ( .IN1(n717), .IN2(n745), .QN(N570) );
  OR2X1 U381 ( .IN1(n899), .IN2(n900), .Q(N57) );
  AO221X1 U382 ( .IN1(n806), .IN2(rdata_1[41]), .IN3(n807), .IN4(rdata_0[41]), 
        .IN5(n901), .Q(n900) );
  AO22X1 U383 ( .IN1(n809), .IN2(rdata_2[41]), .IN3(n720), .IN4(rdata_7[41]), 
        .Q(n901) );
  AO221X1 U384 ( .IN1(n810), .IN2(rdata_4[41]), .IN3(n811), .IN4(rdata_3[41]), 
        .IN5(n902), .Q(n899) );
  AO22X1 U385 ( .IN1(n813), .IN2(rdata_5[41]), .IN3(n814), .IN4(rdata_6[41]), 
        .Q(n902) );
  NOR2X0 U386 ( .IN1(n717), .IN2(n746), .QN(N569) );
  NOR2X0 U387 ( .IN1(n717), .IN2(n747), .QN(N568) );
  NOR2X0 U388 ( .IN1(n717), .IN2(n748), .QN(N567) );
  NOR2X0 U389 ( .IN1(n717), .IN2(n749), .QN(N566) );
  NOR2X0 U390 ( .IN1(n717), .IN2(n750), .QN(N565) );
  NOR2X0 U391 ( .IN1(n717), .IN2(n751), .QN(N564) );
  NOR2X0 U392 ( .IN1(n717), .IN2(n752), .QN(N563) );
  NOR2X0 U393 ( .IN1(n717), .IN2(n753), .QN(N562) );
  NOR2X0 U394 ( .IN1(n717), .IN2(n754), .QN(N561) );
  NOR2X0 U395 ( .IN1(n717), .IN2(n755), .QN(N560) );
  OR2X1 U396 ( .IN1(n903), .IN2(n904), .Q(N56) );
  AO221X1 U397 ( .IN1(n806), .IN2(rdata_1[40]), .IN3(n807), .IN4(rdata_0[40]), 
        .IN5(n905), .Q(n904) );
  AO22X1 U398 ( .IN1(n809), .IN2(rdata_2[40]), .IN3(n720), .IN4(rdata_7[40]), 
        .Q(n905) );
  AO221X1 U399 ( .IN1(n810), .IN2(rdata_4[40]), .IN3(n811), .IN4(rdata_3[40]), 
        .IN5(n906), .Q(n903) );
  AO22X1 U400 ( .IN1(n813), .IN2(rdata_5[40]), .IN3(n814), .IN4(rdata_6[40]), 
        .Q(n906) );
  NOR2X0 U401 ( .IN1(n717), .IN2(n756), .QN(N559) );
  NOR2X0 U402 ( .IN1(n717), .IN2(n757), .QN(N558) );
  NOR2X0 U403 ( .IN1(n717), .IN2(n758), .QN(N557) );
  NOR2X0 U404 ( .IN1(n717), .IN2(n759), .QN(N556) );
  NOR2X0 U405 ( .IN1(n717), .IN2(n760), .QN(N555) );
  NOR2X0 U406 ( .IN1(n717), .IN2(n761), .QN(N554) );
  NOR2X0 U407 ( .IN1(n717), .IN2(n762), .QN(N553) );
  NOR2X0 U408 ( .IN1(n717), .IN2(n763), .QN(N552) );
  NOR2X0 U409 ( .IN1(n717), .IN2(n764), .QN(N551) );
  NOR2X0 U410 ( .IN1(n717), .IN2(n765), .QN(N550) );
  OR2X1 U411 ( .IN1(n907), .IN2(n908), .Q(N55) );
  AO221X1 U412 ( .IN1(n806), .IN2(rdata_1[39]), .IN3(n807), .IN4(rdata_0[39]), 
        .IN5(n909), .Q(n908) );
  AO22X1 U413 ( .IN1(n809), .IN2(rdata_2[39]), .IN3(n720), .IN4(rdata_7[39]), 
        .Q(n909) );
  AO221X1 U414 ( .IN1(n810), .IN2(rdata_4[39]), .IN3(n811), .IN4(rdata_3[39]), 
        .IN5(n910), .Q(n907) );
  AO22X1 U415 ( .IN1(n813), .IN2(rdata_5[39]), .IN3(n814), .IN4(rdata_6[39]), 
        .Q(n910) );
  NOR2X0 U416 ( .IN1(n717), .IN2(n766), .QN(N549) );
  NOR2X0 U417 ( .IN1(n717), .IN2(n767), .QN(N548) );
  NOR2X0 U418 ( .IN1(n717), .IN2(n768), .QN(N547) );
  NOR2X0 U419 ( .IN1(n717), .IN2(n769), .QN(N546) );
  NOR2X0 U420 ( .IN1(n717), .IN2(n770), .QN(N545) );
  NOR2X0 U421 ( .IN1(n717), .IN2(n771), .QN(N544) );
  NOR2X0 U422 ( .IN1(n717), .IN2(n772), .QN(N543) );
  NOR2X0 U423 ( .IN1(n717), .IN2(n773), .QN(N542) );
  NOR2X0 U424 ( .IN1(n717), .IN2(n774), .QN(N541) );
  NOR2X0 U425 ( .IN1(n717), .IN2(n775), .QN(N540) );
  OR2X1 U426 ( .IN1(n911), .IN2(n912), .Q(N54) );
  AO221X1 U427 ( .IN1(n806), .IN2(rdata_1[38]), .IN3(n807), .IN4(rdata_0[38]), 
        .IN5(n913), .Q(n912) );
  AO22X1 U428 ( .IN1(n809), .IN2(rdata_2[38]), .IN3(n720), .IN4(rdata_7[38]), 
        .Q(n913) );
  AO221X1 U429 ( .IN1(n810), .IN2(rdata_4[38]), .IN3(n811), .IN4(rdata_3[38]), 
        .IN5(n914), .Q(n911) );
  AO22X1 U430 ( .IN1(n813), .IN2(rdata_5[38]), .IN3(n814), .IN4(rdata_6[38]), 
        .Q(n914) );
  NOR2X0 U431 ( .IN1(n717), .IN2(n776), .QN(N539) );
  NOR2X0 U432 ( .IN1(n717), .IN2(n777), .QN(N538) );
  NOR2X0 U433 ( .IN1(n717), .IN2(n778), .QN(N537) );
  NOR2X0 U434 ( .IN1(n717), .IN2(n779), .QN(N536) );
  NOR2X0 U435 ( .IN1(n717), .IN2(n780), .QN(N535) );
  NOR2X0 U436 ( .IN1(n717), .IN2(n781), .QN(N534) );
  NOR2X0 U437 ( .IN1(n717), .IN2(n782), .QN(N533) );
  NOR2X0 U438 ( .IN1(n717), .IN2(n783), .QN(N532) );
  NOR2X0 U439 ( .IN1(n717), .IN2(n784), .QN(N531) );
  NOR2X0 U440 ( .IN1(n717), .IN2(n785), .QN(N530) );
  OR2X1 U441 ( .IN1(n915), .IN2(n916), .Q(N53) );
  AO221X1 U442 ( .IN1(n806), .IN2(rdata_1[37]), .IN3(n807), .IN4(rdata_0[37]), 
        .IN5(n917), .Q(n916) );
  AO22X1 U443 ( .IN1(n809), .IN2(rdata_2[37]), .IN3(n720), .IN4(rdata_7[37]), 
        .Q(n917) );
  AO221X1 U444 ( .IN1(n810), .IN2(rdata_4[37]), .IN3(n811), .IN4(rdata_3[37]), 
        .IN5(n918), .Q(n915) );
  AO22X1 U445 ( .IN1(n813), .IN2(rdata_5[37]), .IN3(n814), .IN4(rdata_6[37]), 
        .Q(n918) );
  NOR2X0 U446 ( .IN1(n717), .IN2(n786), .QN(N529) );
  NOR2X0 U447 ( .IN1(n715), .IN2(n723), .QN(N528) );
  NOR2X0 U448 ( .IN1(n715), .IN2(n724), .QN(N527) );
  NOR2X0 U449 ( .IN1(n715), .IN2(n725), .QN(N526) );
  NOR2X0 U450 ( .IN1(n715), .IN2(n726), .QN(N525) );
  NOR2X0 U451 ( .IN1(n715), .IN2(n727), .QN(N524) );
  NOR2X0 U452 ( .IN1(n715), .IN2(n728), .QN(N523) );
  NOR2X0 U453 ( .IN1(n715), .IN2(n729), .QN(N522) );
  NOR2X0 U454 ( .IN1(n715), .IN2(n730), .QN(N521) );
  NOR2X0 U455 ( .IN1(n715), .IN2(n731), .QN(N520) );
  OR2X1 U456 ( .IN1(n919), .IN2(n920), .Q(N52) );
  AO221X1 U457 ( .IN1(n806), .IN2(rdata_1[36]), .IN3(n807), .IN4(rdata_0[36]), 
        .IN5(n921), .Q(n920) );
  AO22X1 U458 ( .IN1(n809), .IN2(rdata_2[36]), .IN3(n720), .IN4(rdata_7[36]), 
        .Q(n921) );
  AO221X1 U459 ( .IN1(n810), .IN2(rdata_4[36]), .IN3(n811), .IN4(rdata_3[36]), 
        .IN5(n922), .Q(n919) );
  AO22X1 U460 ( .IN1(n813), .IN2(rdata_5[36]), .IN3(n814), .IN4(rdata_6[36]), 
        .Q(n922) );
  NOR2X0 U461 ( .IN1(n715), .IN2(n732), .QN(N519) );
  NOR2X0 U462 ( .IN1(n715), .IN2(n733), .QN(N518) );
  NOR2X0 U463 ( .IN1(n715), .IN2(n734), .QN(N517) );
  NOR2X0 U464 ( .IN1(n715), .IN2(n735), .QN(N516) );
  NOR2X0 U465 ( .IN1(n715), .IN2(n736), .QN(N515) );
  NOR2X0 U466 ( .IN1(n715), .IN2(n737), .QN(N514) );
  NOR2X0 U467 ( .IN1(n715), .IN2(n738), .QN(N513) );
  NOR2X0 U468 ( .IN1(n715), .IN2(n739), .QN(N512) );
  NOR2X0 U469 ( .IN1(n715), .IN2(n740), .QN(N511) );
  NOR2X0 U470 ( .IN1(n715), .IN2(n741), .QN(N510) );
  OR2X1 U471 ( .IN1(n923), .IN2(n924), .Q(N51) );
  AO221X1 U472 ( .IN1(n806), .IN2(rdata_1[35]), .IN3(n807), .IN4(rdata_0[35]), 
        .IN5(n925), .Q(n924) );
  AO22X1 U473 ( .IN1(n809), .IN2(rdata_2[35]), .IN3(n720), .IN4(rdata_7[35]), 
        .Q(n925) );
  AO221X1 U474 ( .IN1(n810), .IN2(rdata_4[35]), .IN3(n811), .IN4(rdata_3[35]), 
        .IN5(n926), .Q(n923) );
  AO22X1 U475 ( .IN1(n813), .IN2(rdata_5[35]), .IN3(n814), .IN4(rdata_6[35]), 
        .Q(n926) );
  NOR2X0 U476 ( .IN1(n715), .IN2(n742), .QN(N509) );
  NOR2X0 U477 ( .IN1(n715), .IN2(n743), .QN(N508) );
  NOR2X0 U478 ( .IN1(n715), .IN2(n744), .QN(N507) );
  NOR2X0 U479 ( .IN1(n715), .IN2(n745), .QN(N506) );
  NOR2X0 U480 ( .IN1(n715), .IN2(n746), .QN(N505) );
  NOR2X0 U481 ( .IN1(n715), .IN2(n747), .QN(N504) );
  NOR2X0 U482 ( .IN1(n715), .IN2(n748), .QN(N503) );
  NOR2X0 U483 ( .IN1(n715), .IN2(n749), .QN(N502) );
  NOR2X0 U484 ( .IN1(n715), .IN2(n750), .QN(N501) );
  NOR2X0 U485 ( .IN1(n715), .IN2(n751), .QN(N500) );
  OR2X1 U486 ( .IN1(n927), .IN2(n928), .Q(N50) );
  AO221X1 U487 ( .IN1(n806), .IN2(rdata_1[34]), .IN3(n807), .IN4(rdata_0[34]), 
        .IN5(n929), .Q(n928) );
  AO22X1 U488 ( .IN1(n809), .IN2(rdata_2[34]), .IN3(n720), .IN4(rdata_7[34]), 
        .Q(n929) );
  AO221X1 U489 ( .IN1(n810), .IN2(rdata_4[34]), .IN3(n811), .IN4(rdata_3[34]), 
        .IN5(n930), .Q(n927) );
  AO22X1 U490 ( .IN1(n813), .IN2(rdata_5[34]), .IN3(n814), .IN4(rdata_6[34]), 
        .Q(n930) );
  NOR2X0 U491 ( .IN1(n715), .IN2(n752), .QN(N499) );
  NOR2X0 U492 ( .IN1(n715), .IN2(n753), .QN(N498) );
  NOR2X0 U493 ( .IN1(n715), .IN2(n754), .QN(N497) );
  NOR2X0 U494 ( .IN1(n715), .IN2(n755), .QN(N496) );
  NOR2X0 U495 ( .IN1(n715), .IN2(n756), .QN(N495) );
  NOR2X0 U496 ( .IN1(n715), .IN2(n757), .QN(N494) );
  NOR2X0 U497 ( .IN1(n715), .IN2(n758), .QN(N493) );
  NOR2X0 U498 ( .IN1(n715), .IN2(n759), .QN(N492) );
  NOR2X0 U499 ( .IN1(n715), .IN2(n760), .QN(N491) );
  NOR2X0 U500 ( .IN1(n715), .IN2(n761), .QN(N490) );
  OR2X1 U501 ( .IN1(n931), .IN2(n932), .Q(N49) );
  AO221X1 U502 ( .IN1(n806), .IN2(rdata_1[33]), .IN3(n807), .IN4(rdata_0[33]), 
        .IN5(n933), .Q(n932) );
  AO22X1 U503 ( .IN1(n809), .IN2(rdata_2[33]), .IN3(n720), .IN4(rdata_7[33]), 
        .Q(n933) );
  AO221X1 U504 ( .IN1(n810), .IN2(rdata_4[33]), .IN3(n811), .IN4(rdata_3[33]), 
        .IN5(n934), .Q(n931) );
  AO22X1 U505 ( .IN1(n813), .IN2(rdata_5[33]), .IN3(n814), .IN4(rdata_6[33]), 
        .Q(n934) );
  NOR2X0 U506 ( .IN1(n715), .IN2(n762), .QN(N489) );
  NOR2X0 U507 ( .IN1(n715), .IN2(n763), .QN(N488) );
  NOR2X0 U508 ( .IN1(n715), .IN2(n764), .QN(N487) );
  NOR2X0 U509 ( .IN1(n715), .IN2(n765), .QN(N486) );
  NOR2X0 U510 ( .IN1(n715), .IN2(n766), .QN(N485) );
  NOR2X0 U511 ( .IN1(n715), .IN2(n767), .QN(N484) );
  NOR2X0 U512 ( .IN1(n715), .IN2(n768), .QN(N483) );
  NOR2X0 U513 ( .IN1(n715), .IN2(n769), .QN(N482) );
  NOR2X0 U514 ( .IN1(n715), .IN2(n770), .QN(N481) );
  NOR2X0 U515 ( .IN1(n715), .IN2(n771), .QN(N480) );
  OR2X1 U516 ( .IN1(n935), .IN2(n936), .Q(N48) );
  AO221X1 U517 ( .IN1(n806), .IN2(rdata_1[32]), .IN3(n807), .IN4(rdata_0[32]), 
        .IN5(n937), .Q(n936) );
  AO22X1 U518 ( .IN1(n809), .IN2(rdata_2[32]), .IN3(n720), .IN4(rdata_7[32]), 
        .Q(n937) );
  AO221X1 U519 ( .IN1(n810), .IN2(rdata_4[32]), .IN3(n811), .IN4(rdata_3[32]), 
        .IN5(n938), .Q(n935) );
  AO22X1 U520 ( .IN1(n813), .IN2(rdata_5[32]), .IN3(n814), .IN4(rdata_6[32]), 
        .Q(n938) );
  NOR2X0 U521 ( .IN1(n715), .IN2(n772), .QN(N479) );
  NOR2X0 U522 ( .IN1(n715), .IN2(n773), .QN(N478) );
  NOR2X0 U523 ( .IN1(n715), .IN2(n774), .QN(N477) );
  NOR2X0 U524 ( .IN1(n715), .IN2(n775), .QN(N476) );
  NOR2X0 U525 ( .IN1(n715), .IN2(n776), .QN(N475) );
  NOR2X0 U526 ( .IN1(n715), .IN2(n777), .QN(N474) );
  NOR2X0 U527 ( .IN1(n715), .IN2(n778), .QN(N473) );
  NOR2X0 U528 ( .IN1(n715), .IN2(n779), .QN(N472) );
  NOR2X0 U529 ( .IN1(n715), .IN2(n780), .QN(N471) );
  NOR2X0 U530 ( .IN1(n715), .IN2(n781), .QN(N470) );
  OR2X1 U531 ( .IN1(n939), .IN2(n940), .Q(N47) );
  AO221X1 U532 ( .IN1(n806), .IN2(rdata_1[31]), .IN3(n807), .IN4(rdata_0[31]), 
        .IN5(n941), .Q(n940) );
  AO22X1 U533 ( .IN1(n809), .IN2(rdata_2[31]), .IN3(n720), .IN4(rdata_7[31]), 
        .Q(n941) );
  AO221X1 U534 ( .IN1(n810), .IN2(rdata_4[31]), .IN3(n811), .IN4(rdata_3[31]), 
        .IN5(n942), .Q(n939) );
  AO22X1 U535 ( .IN1(n813), .IN2(rdata_5[31]), .IN3(n814), .IN4(rdata_6[31]), 
        .Q(n942) );
  NOR2X0 U536 ( .IN1(n715), .IN2(n782), .QN(N469) );
  NOR2X0 U537 ( .IN1(n715), .IN2(n783), .QN(N468) );
  NOR2X0 U538 ( .IN1(n715), .IN2(n784), .QN(N467) );
  NOR2X0 U539 ( .IN1(n715), .IN2(n785), .QN(N466) );
  NOR2X0 U540 ( .IN1(n715), .IN2(n786), .QN(N465) );
  NOR2X0 U541 ( .IN1(n716), .IN2(n723), .QN(N464) );
  NOR2X0 U542 ( .IN1(n716), .IN2(n724), .QN(N463) );
  NOR2X0 U543 ( .IN1(n716), .IN2(n725), .QN(N462) );
  NOR2X0 U544 ( .IN1(n716), .IN2(n726), .QN(N461) );
  NOR2X0 U545 ( .IN1(n716), .IN2(n727), .QN(N460) );
  OR2X1 U546 ( .IN1(n943), .IN2(n944), .Q(N46) );
  AO221X1 U547 ( .IN1(n806), .IN2(rdata_1[30]), .IN3(n807), .IN4(rdata_0[30]), 
        .IN5(n945), .Q(n944) );
  AO22X1 U548 ( .IN1(n809), .IN2(rdata_2[30]), .IN3(n720), .IN4(rdata_7[30]), 
        .Q(n945) );
  AO221X1 U549 ( .IN1(n810), .IN2(rdata_4[30]), .IN3(n811), .IN4(rdata_3[30]), 
        .IN5(n946), .Q(n943) );
  AO22X1 U550 ( .IN1(n813), .IN2(rdata_5[30]), .IN3(n814), .IN4(rdata_6[30]), 
        .Q(n946) );
  NOR2X0 U551 ( .IN1(n716), .IN2(n728), .QN(N459) );
  NOR2X0 U552 ( .IN1(n716), .IN2(n729), .QN(N458) );
  NOR2X0 U553 ( .IN1(n716), .IN2(n730), .QN(N457) );
  NOR2X0 U554 ( .IN1(n716), .IN2(n731), .QN(N456) );
  NOR2X0 U555 ( .IN1(n716), .IN2(n732), .QN(N455) );
  NOR2X0 U556 ( .IN1(n716), .IN2(n733), .QN(N454) );
  NOR2X0 U557 ( .IN1(n716), .IN2(n734), .QN(N453) );
  NOR2X0 U558 ( .IN1(n716), .IN2(n735), .QN(N452) );
  NOR2X0 U559 ( .IN1(n716), .IN2(n736), .QN(N451) );
  NOR2X0 U560 ( .IN1(n716), .IN2(n737), .QN(N450) );
  OR2X1 U561 ( .IN1(n947), .IN2(n948), .Q(N45) );
  AO221X1 U562 ( .IN1(n806), .IN2(rdata_1[29]), .IN3(n807), .IN4(rdata_0[29]), 
        .IN5(n949), .Q(n948) );
  AO22X1 U563 ( .IN1(n809), .IN2(rdata_2[29]), .IN3(n720), .IN4(rdata_7[29]), 
        .Q(n949) );
  AO221X1 U564 ( .IN1(n810), .IN2(rdata_4[29]), .IN3(n811), .IN4(rdata_3[29]), 
        .IN5(n950), .Q(n947) );
  AO22X1 U565 ( .IN1(n813), .IN2(rdata_5[29]), .IN3(n814), .IN4(rdata_6[29]), 
        .Q(n950) );
  NOR2X0 U566 ( .IN1(n716), .IN2(n738), .QN(N449) );
  NOR2X0 U567 ( .IN1(n716), .IN2(n739), .QN(N448) );
  NOR2X0 U568 ( .IN1(n716), .IN2(n740), .QN(N447) );
  NOR2X0 U569 ( .IN1(n716), .IN2(n741), .QN(N446) );
  NOR2X0 U570 ( .IN1(n716), .IN2(n742), .QN(N445) );
  NOR2X0 U571 ( .IN1(n716), .IN2(n743), .QN(N444) );
  NOR2X0 U572 ( .IN1(n716), .IN2(n744), .QN(N443) );
  NOR2X0 U573 ( .IN1(n716), .IN2(n745), .QN(N442) );
  NOR2X0 U574 ( .IN1(n716), .IN2(n746), .QN(N441) );
  NOR2X0 U575 ( .IN1(n716), .IN2(n747), .QN(N440) );
  OR2X1 U576 ( .IN1(n951), .IN2(n952), .Q(N44) );
  AO221X1 U577 ( .IN1(n806), .IN2(rdata_1[28]), .IN3(n807), .IN4(rdata_0[28]), 
        .IN5(n953), .Q(n952) );
  AO22X1 U578 ( .IN1(n809), .IN2(rdata_2[28]), .IN3(n720), .IN4(rdata_7[28]), 
        .Q(n953) );
  AO221X1 U579 ( .IN1(n810), .IN2(rdata_4[28]), .IN3(n811), .IN4(rdata_3[28]), 
        .IN5(n954), .Q(n951) );
  AO22X1 U580 ( .IN1(n813), .IN2(rdata_5[28]), .IN3(n814), .IN4(rdata_6[28]), 
        .Q(n954) );
  NOR2X0 U581 ( .IN1(n716), .IN2(n748), .QN(N439) );
  NOR2X0 U582 ( .IN1(n716), .IN2(n749), .QN(N438) );
  NOR2X0 U583 ( .IN1(n716), .IN2(n750), .QN(N437) );
  NOR2X0 U584 ( .IN1(n716), .IN2(n751), .QN(N436) );
  NOR2X0 U585 ( .IN1(n716), .IN2(n752), .QN(N435) );
  NOR2X0 U586 ( .IN1(n716), .IN2(n753), .QN(N434) );
  NOR2X0 U587 ( .IN1(n716), .IN2(n754), .QN(N433) );
  NOR2X0 U588 ( .IN1(n716), .IN2(n755), .QN(N432) );
  NOR2X0 U589 ( .IN1(n716), .IN2(n756), .QN(N431) );
  NOR2X0 U590 ( .IN1(n716), .IN2(n757), .QN(N430) );
  OR2X1 U591 ( .IN1(n955), .IN2(n956), .Q(N43) );
  AO221X1 U592 ( .IN1(n806), .IN2(rdata_1[27]), .IN3(n807), .IN4(rdata_0[27]), 
        .IN5(n957), .Q(n956) );
  AO22X1 U593 ( .IN1(n809), .IN2(rdata_2[27]), .IN3(n720), .IN4(rdata_7[27]), 
        .Q(n957) );
  AO221X1 U594 ( .IN1(n810), .IN2(rdata_4[27]), .IN3(n811), .IN4(rdata_3[27]), 
        .IN5(n958), .Q(n955) );
  AO22X1 U595 ( .IN1(n813), .IN2(rdata_5[27]), .IN3(n814), .IN4(rdata_6[27]), 
        .Q(n958) );
  NOR2X0 U596 ( .IN1(n716), .IN2(n758), .QN(N429) );
  NOR2X0 U597 ( .IN1(n716), .IN2(n759), .QN(N428) );
  NOR2X0 U598 ( .IN1(n716), .IN2(n760), .QN(N427) );
  NOR2X0 U599 ( .IN1(n716), .IN2(n761), .QN(N426) );
  NOR2X0 U600 ( .IN1(n716), .IN2(n762), .QN(N425) );
  NOR2X0 U601 ( .IN1(n716), .IN2(n763), .QN(N424) );
  NOR2X0 U602 ( .IN1(n716), .IN2(n764), .QN(N423) );
  NOR2X0 U603 ( .IN1(n716), .IN2(n765), .QN(N422) );
  NOR2X0 U604 ( .IN1(n716), .IN2(n766), .QN(N421) );
  NOR2X0 U605 ( .IN1(n716), .IN2(n767), .QN(N420) );
  OR2X1 U606 ( .IN1(n959), .IN2(n960), .Q(N42) );
  AO221X1 U607 ( .IN1(n806), .IN2(rdata_1[26]), .IN3(n807), .IN4(rdata_0[26]), 
        .IN5(n961), .Q(n960) );
  AO22X1 U608 ( .IN1(n809), .IN2(rdata_2[26]), .IN3(n720), .IN4(rdata_7[26]), 
        .Q(n961) );
  AO221X1 U609 ( .IN1(n810), .IN2(rdata_4[26]), .IN3(n811), .IN4(rdata_3[26]), 
        .IN5(n962), .Q(n959) );
  AO22X1 U610 ( .IN1(n813), .IN2(rdata_5[26]), .IN3(n814), .IN4(rdata_6[26]), 
        .Q(n962) );
  NOR2X0 U611 ( .IN1(n716), .IN2(n768), .QN(N419) );
  NOR2X0 U612 ( .IN1(n716), .IN2(n769), .QN(N418) );
  NOR2X0 U613 ( .IN1(n716), .IN2(n770), .QN(N417) );
  NOR2X0 U614 ( .IN1(n716), .IN2(n771), .QN(N416) );
  NOR2X0 U615 ( .IN1(n716), .IN2(n772), .QN(N415) );
  NOR2X0 U616 ( .IN1(n716), .IN2(n773), .QN(N414) );
  NOR2X0 U617 ( .IN1(n716), .IN2(n774), .QN(N413) );
  NOR2X0 U618 ( .IN1(n716), .IN2(n775), .QN(N412) );
  NOR2X0 U619 ( .IN1(n716), .IN2(n776), .QN(N411) );
  NOR2X0 U620 ( .IN1(n716), .IN2(n777), .QN(N410) );
  OR2X1 U621 ( .IN1(n963), .IN2(n964), .Q(N41) );
  AO221X1 U622 ( .IN1(n806), .IN2(rdata_1[25]), .IN3(n807), .IN4(rdata_0[25]), 
        .IN5(n965), .Q(n964) );
  AO22X1 U623 ( .IN1(n809), .IN2(rdata_2[25]), .IN3(n720), .IN4(rdata_7[25]), 
        .Q(n965) );
  AO221X1 U624 ( .IN1(n810), .IN2(rdata_4[25]), .IN3(n811), .IN4(rdata_3[25]), 
        .IN5(n966), .Q(n963) );
  AO22X1 U625 ( .IN1(n813), .IN2(rdata_5[25]), .IN3(n814), .IN4(rdata_6[25]), 
        .Q(n966) );
  NOR2X0 U626 ( .IN1(n716), .IN2(n778), .QN(N409) );
  NOR2X0 U627 ( .IN1(n716), .IN2(n779), .QN(N408) );
  NOR2X0 U628 ( .IN1(n716), .IN2(n780), .QN(N407) );
  NOR2X0 U629 ( .IN1(n716), .IN2(n781), .QN(N406) );
  NOR2X0 U630 ( .IN1(n716), .IN2(n782), .QN(N405) );
  NOR2X0 U631 ( .IN1(n716), .IN2(n783), .QN(N404) );
  NOR2X0 U632 ( .IN1(n716), .IN2(n784), .QN(N403) );
  NOR2X0 U633 ( .IN1(n716), .IN2(n785), .QN(N402) );
  NOR2X0 U634 ( .IN1(n716), .IN2(n786), .QN(N401) );
  NOR2X0 U635 ( .IN1(n714), .IN2(n723), .QN(N400) );
  OR2X1 U636 ( .IN1(n967), .IN2(n968), .Q(N40) );
  AO221X1 U637 ( .IN1(n806), .IN2(rdata_1[24]), .IN3(n807), .IN4(rdata_0[24]), 
        .IN5(n969), .Q(n968) );
  AO22X1 U638 ( .IN1(n809), .IN2(rdata_2[24]), .IN3(n720), .IN4(rdata_7[24]), 
        .Q(n969) );
  AO221X1 U639 ( .IN1(n810), .IN2(rdata_4[24]), .IN3(n811), .IN4(rdata_3[24]), 
        .IN5(n970), .Q(n967) );
  AO22X1 U640 ( .IN1(n813), .IN2(rdata_5[24]), .IN3(n814), .IN4(rdata_6[24]), 
        .Q(n970) );
  NOR2X0 U641 ( .IN1(n714), .IN2(n724), .QN(N399) );
  NOR2X0 U642 ( .IN1(n714), .IN2(n725), .QN(N398) );
  NOR2X0 U643 ( .IN1(n714), .IN2(n726), .QN(N397) );
  NOR2X0 U644 ( .IN1(n714), .IN2(n727), .QN(N396) );
  NOR2X0 U645 ( .IN1(n714), .IN2(n728), .QN(N395) );
  NOR2X0 U646 ( .IN1(n714), .IN2(n729), .QN(N394) );
  NOR2X0 U647 ( .IN1(n714), .IN2(n730), .QN(N393) );
  NOR2X0 U648 ( .IN1(n714), .IN2(n731), .QN(N392) );
  NOR2X0 U649 ( .IN1(n714), .IN2(n732), .QN(N391) );
  NOR2X0 U650 ( .IN1(n714), .IN2(n733), .QN(N390) );
  OR2X1 U651 ( .IN1(n971), .IN2(n972), .Q(N39) );
  AO221X1 U652 ( .IN1(n806), .IN2(rdata_1[23]), .IN3(n807), .IN4(rdata_0[23]), 
        .IN5(n973), .Q(n972) );
  AO22X1 U653 ( .IN1(n809), .IN2(rdata_2[23]), .IN3(n720), .IN4(rdata_7[23]), 
        .Q(n973) );
  AO221X1 U654 ( .IN1(n810), .IN2(rdata_4[23]), .IN3(n811), .IN4(rdata_3[23]), 
        .IN5(n974), .Q(n971) );
  AO22X1 U655 ( .IN1(n813), .IN2(rdata_5[23]), .IN3(n814), .IN4(rdata_6[23]), 
        .Q(n974) );
  NOR2X0 U656 ( .IN1(n714), .IN2(n734), .QN(N389) );
  NOR2X0 U657 ( .IN1(n714), .IN2(n735), .QN(N388) );
  NOR2X0 U658 ( .IN1(n714), .IN2(n736), .QN(N387) );
  NOR2X0 U659 ( .IN1(n714), .IN2(n737), .QN(N386) );
  NOR2X0 U660 ( .IN1(n714), .IN2(n738), .QN(N385) );
  NOR2X0 U661 ( .IN1(n714), .IN2(n739), .QN(N384) );
  NOR2X0 U662 ( .IN1(n714), .IN2(n740), .QN(N383) );
  NOR2X0 U663 ( .IN1(n714), .IN2(n741), .QN(N382) );
  NOR2X0 U664 ( .IN1(n714), .IN2(n742), .QN(N381) );
  NOR2X0 U665 ( .IN1(n714), .IN2(n743), .QN(N380) );
  OR2X1 U666 ( .IN1(n975), .IN2(n976), .Q(N38) );
  AO221X1 U667 ( .IN1(n806), .IN2(rdata_1[22]), .IN3(n807), .IN4(rdata_0[22]), 
        .IN5(n977), .Q(n976) );
  AO22X1 U668 ( .IN1(n809), .IN2(rdata_2[22]), .IN3(n720), .IN4(rdata_7[22]), 
        .Q(n977) );
  AO221X1 U669 ( .IN1(n810), .IN2(rdata_4[22]), .IN3(n811), .IN4(rdata_3[22]), 
        .IN5(n978), .Q(n975) );
  AO22X1 U670 ( .IN1(n813), .IN2(rdata_5[22]), .IN3(n814), .IN4(rdata_6[22]), 
        .Q(n978) );
  NOR2X0 U671 ( .IN1(n714), .IN2(n744), .QN(N379) );
  NOR2X0 U672 ( .IN1(n714), .IN2(n745), .QN(N378) );
  NOR2X0 U673 ( .IN1(n714), .IN2(n746), .QN(N377) );
  NOR2X0 U674 ( .IN1(n714), .IN2(n747), .QN(N376) );
  NOR2X0 U675 ( .IN1(n714), .IN2(n748), .QN(N375) );
  NOR2X0 U676 ( .IN1(n714), .IN2(n749), .QN(N374) );
  NOR2X0 U677 ( .IN1(n714), .IN2(n750), .QN(N373) );
  NOR2X0 U678 ( .IN1(n714), .IN2(n751), .QN(N372) );
  NOR2X0 U679 ( .IN1(n714), .IN2(n752), .QN(N371) );
  NOR2X0 U680 ( .IN1(n714), .IN2(n753), .QN(N370) );
  OR2X1 U681 ( .IN1(n979), .IN2(n980), .Q(N37) );
  AO221X1 U682 ( .IN1(n806), .IN2(rdata_1[21]), .IN3(n807), .IN4(rdata_0[21]), 
        .IN5(n981), .Q(n980) );
  AO22X1 U683 ( .IN1(n809), .IN2(rdata_2[21]), .IN3(n720), .IN4(rdata_7[21]), 
        .Q(n981) );
  AO221X1 U684 ( .IN1(n810), .IN2(rdata_4[21]), .IN3(n811), .IN4(rdata_3[21]), 
        .IN5(n982), .Q(n979) );
  AO22X1 U685 ( .IN1(n813), .IN2(rdata_5[21]), .IN3(n814), .IN4(rdata_6[21]), 
        .Q(n982) );
  NOR2X0 U686 ( .IN1(n714), .IN2(n754), .QN(N369) );
  NOR2X0 U687 ( .IN1(n714), .IN2(n755), .QN(N368) );
  NOR2X0 U688 ( .IN1(n714), .IN2(n756), .QN(N367) );
  NOR2X0 U689 ( .IN1(n714), .IN2(n757), .QN(N366) );
  NOR2X0 U690 ( .IN1(n714), .IN2(n758), .QN(N365) );
  NOR2X0 U691 ( .IN1(n714), .IN2(n759), .QN(N364) );
  NOR2X0 U692 ( .IN1(n714), .IN2(n760), .QN(N363) );
  NOR2X0 U693 ( .IN1(n714), .IN2(n761), .QN(N362) );
  NOR2X0 U694 ( .IN1(n714), .IN2(n762), .QN(N361) );
  NOR2X0 U695 ( .IN1(n714), .IN2(n763), .QN(N360) );
  OR2X1 U696 ( .IN1(n983), .IN2(n984), .Q(N36) );
  AO221X1 U697 ( .IN1(n806), .IN2(rdata_1[20]), .IN3(n807), .IN4(rdata_0[20]), 
        .IN5(n985), .Q(n984) );
  AO22X1 U698 ( .IN1(n809), .IN2(rdata_2[20]), .IN3(n720), .IN4(rdata_7[20]), 
        .Q(n985) );
  AO221X1 U699 ( .IN1(n810), .IN2(rdata_4[20]), .IN3(n811), .IN4(rdata_3[20]), 
        .IN5(n986), .Q(n983) );
  AO22X1 U700 ( .IN1(n813), .IN2(rdata_5[20]), .IN3(n814), .IN4(rdata_6[20]), 
        .Q(n986) );
  NOR2X0 U701 ( .IN1(n714), .IN2(n764), .QN(N359) );
  NOR2X0 U702 ( .IN1(n714), .IN2(n765), .QN(N358) );
  NOR2X0 U703 ( .IN1(n714), .IN2(n766), .QN(N357) );
  NOR2X0 U704 ( .IN1(n714), .IN2(n767), .QN(N356) );
  NOR2X0 U705 ( .IN1(n714), .IN2(n768), .QN(N355) );
  NOR2X0 U706 ( .IN1(n714), .IN2(n769), .QN(N354) );
  NOR2X0 U707 ( .IN1(n714), .IN2(n770), .QN(N353) );
  NOR2X0 U708 ( .IN1(n714), .IN2(n771), .QN(N352) );
  NOR2X0 U709 ( .IN1(n714), .IN2(n772), .QN(N351) );
  NOR2X0 U710 ( .IN1(n714), .IN2(n773), .QN(N350) );
  OR2X1 U711 ( .IN1(n987), .IN2(n988), .Q(N35) );
  AO221X1 U712 ( .IN1(n806), .IN2(rdata_1[19]), .IN3(n807), .IN4(rdata_0[19]), 
        .IN5(n989), .Q(n988) );
  AO22X1 U713 ( .IN1(n809), .IN2(rdata_2[19]), .IN3(n720), .IN4(rdata_7[19]), 
        .Q(n989) );
  AO221X1 U714 ( .IN1(n810), .IN2(rdata_4[19]), .IN3(n811), .IN4(rdata_3[19]), 
        .IN5(n990), .Q(n987) );
  AO22X1 U715 ( .IN1(n813), .IN2(rdata_5[19]), .IN3(n814), .IN4(rdata_6[19]), 
        .Q(n990) );
  NOR2X0 U716 ( .IN1(n714), .IN2(n774), .QN(N349) );
  NOR2X0 U717 ( .IN1(n714), .IN2(n775), .QN(N348) );
  NOR2X0 U718 ( .IN1(n714), .IN2(n776), .QN(N347) );
  NOR2X0 U719 ( .IN1(n714), .IN2(n777), .QN(N346) );
  NOR2X0 U720 ( .IN1(n714), .IN2(n778), .QN(N345) );
  NOR2X0 U721 ( .IN1(n714), .IN2(n779), .QN(N344) );
  NOR2X0 U722 ( .IN1(n714), .IN2(n780), .QN(N343) );
  NOR2X0 U723 ( .IN1(n714), .IN2(n781), .QN(N342) );
  NOR2X0 U724 ( .IN1(n714), .IN2(n782), .QN(N341) );
  NOR2X0 U725 ( .IN1(n714), .IN2(n783), .QN(N340) );
  OR2X1 U726 ( .IN1(n991), .IN2(n992), .Q(N34) );
  AO221X1 U727 ( .IN1(n806), .IN2(rdata_1[18]), .IN3(n807), .IN4(rdata_0[18]), 
        .IN5(n993), .Q(n992) );
  AO22X1 U728 ( .IN1(n809), .IN2(rdata_2[18]), .IN3(n720), .IN4(rdata_7[18]), 
        .Q(n993) );
  AO221X1 U729 ( .IN1(n810), .IN2(rdata_4[18]), .IN3(n811), .IN4(rdata_3[18]), 
        .IN5(n994), .Q(n991) );
  AO22X1 U730 ( .IN1(n813), .IN2(rdata_5[18]), .IN3(n814), .IN4(rdata_6[18]), 
        .Q(n994) );
  NOR2X0 U731 ( .IN1(n714), .IN2(n784), .QN(N339) );
  NOR2X0 U732 ( .IN1(n714), .IN2(n785), .QN(N338) );
  NOR2X0 U733 ( .IN1(n714), .IN2(n786), .QN(N337) );
  NOR2X0 U734 ( .IN1(n713), .IN2(n723), .QN(N336) );
  NOR2X0 U735 ( .IN1(n713), .IN2(n724), .QN(N335) );
  NOR2X0 U736 ( .IN1(n713), .IN2(n725), .QN(N334) );
  NOR2X0 U737 ( .IN1(n713), .IN2(n726), .QN(N333) );
  NOR2X0 U738 ( .IN1(n713), .IN2(n727), .QN(N332) );
  NOR2X0 U739 ( .IN1(n713), .IN2(n728), .QN(N331) );
  NOR2X0 U740 ( .IN1(n713), .IN2(n729), .QN(N330) );
  OR2X1 U741 ( .IN1(n995), .IN2(n996), .Q(N33) );
  AO221X1 U742 ( .IN1(n806), .IN2(rdata_1[17]), .IN3(n807), .IN4(rdata_0[17]), 
        .IN5(n997), .Q(n996) );
  AO22X1 U743 ( .IN1(n809), .IN2(rdata_2[17]), .IN3(n720), .IN4(rdata_7[17]), 
        .Q(n997) );
  AO221X1 U744 ( .IN1(n810), .IN2(rdata_4[17]), .IN3(n811), .IN4(rdata_3[17]), 
        .IN5(n998), .Q(n995) );
  AO22X1 U745 ( .IN1(n813), .IN2(rdata_5[17]), .IN3(n814), .IN4(rdata_6[17]), 
        .Q(n998) );
  NOR2X0 U746 ( .IN1(n713), .IN2(n730), .QN(N329) );
  NOR2X0 U747 ( .IN1(n713), .IN2(n731), .QN(N328) );
  NOR2X0 U748 ( .IN1(n713), .IN2(n732), .QN(N327) );
  NOR2X0 U749 ( .IN1(n713), .IN2(n733), .QN(N326) );
  NOR2X0 U750 ( .IN1(n713), .IN2(n734), .QN(N325) );
  NOR2X0 U751 ( .IN1(n713), .IN2(n735), .QN(N324) );
  NOR2X0 U752 ( .IN1(n713), .IN2(n736), .QN(N323) );
  NOR2X0 U753 ( .IN1(n713), .IN2(n737), .QN(N322) );
  NOR2X0 U754 ( .IN1(n713), .IN2(n738), .QN(N321) );
  NOR2X0 U755 ( .IN1(n713), .IN2(n739), .QN(N320) );
  OR2X1 U756 ( .IN1(n999), .IN2(n1000), .Q(N32) );
  AO221X1 U757 ( .IN1(n806), .IN2(rdata_1[16]), .IN3(n807), .IN4(rdata_0[16]), 
        .IN5(n1001), .Q(n1000) );
  AO22X1 U758 ( .IN1(n809), .IN2(rdata_2[16]), .IN3(n720), .IN4(rdata_7[16]), 
        .Q(n1001) );
  AO221X1 U759 ( .IN1(n810), .IN2(rdata_4[16]), .IN3(n811), .IN4(rdata_3[16]), 
        .IN5(n1002), .Q(n999) );
  AO22X1 U760 ( .IN1(n813), .IN2(rdata_5[16]), .IN3(n814), .IN4(rdata_6[16]), 
        .Q(n1002) );
  NOR2X0 U761 ( .IN1(n713), .IN2(n740), .QN(N319) );
  NOR2X0 U762 ( .IN1(n713), .IN2(n741), .QN(N318) );
  NOR2X0 U763 ( .IN1(n713), .IN2(n742), .QN(N317) );
  NOR2X0 U764 ( .IN1(n713), .IN2(n743), .QN(N316) );
  NOR2X0 U765 ( .IN1(n713), .IN2(n744), .QN(N315) );
  NOR2X0 U766 ( .IN1(n713), .IN2(n745), .QN(N314) );
  NOR2X0 U767 ( .IN1(n713), .IN2(n746), .QN(N313) );
  NOR2X0 U768 ( .IN1(n713), .IN2(n747), .QN(N312) );
  NOR2X0 U769 ( .IN1(n713), .IN2(n748), .QN(N311) );
  NOR2X0 U770 ( .IN1(n713), .IN2(n749), .QN(N310) );
  OR2X1 U771 ( .IN1(n1003), .IN2(n1004), .Q(N31) );
  AO221X1 U772 ( .IN1(n806), .IN2(rdata_1[15]), .IN3(n807), .IN4(rdata_0[15]), 
        .IN5(n1005), .Q(n1004) );
  AO22X1 U773 ( .IN1(n809), .IN2(rdata_2[15]), .IN3(n720), .IN4(rdata_7[15]), 
        .Q(n1005) );
  AO221X1 U774 ( .IN1(n810), .IN2(rdata_4[15]), .IN3(n811), .IN4(rdata_3[15]), 
        .IN5(n1006), .Q(n1003) );
  AO22X1 U775 ( .IN1(n813), .IN2(rdata_5[15]), .IN3(n814), .IN4(rdata_6[15]), 
        .Q(n1006) );
  NOR2X0 U776 ( .IN1(n713), .IN2(n750), .QN(N309) );
  NOR2X0 U777 ( .IN1(n713), .IN2(n751), .QN(N308) );
  NOR2X0 U778 ( .IN1(n713), .IN2(n752), .QN(N307) );
  NOR2X0 U779 ( .IN1(n713), .IN2(n753), .QN(N306) );
  NOR2X0 U780 ( .IN1(n713), .IN2(n754), .QN(N305) );
  NOR2X0 U781 ( .IN1(n713), .IN2(n755), .QN(N304) );
  NOR2X0 U782 ( .IN1(n713), .IN2(n756), .QN(N303) );
  NOR2X0 U783 ( .IN1(n713), .IN2(n757), .QN(N302) );
  NOR2X0 U784 ( .IN1(n713), .IN2(n758), .QN(N301) );
  NOR2X0 U785 ( .IN1(n713), .IN2(n759), .QN(N300) );
  OR2X1 U786 ( .IN1(n1007), .IN2(n1008), .Q(N30) );
  AO221X1 U787 ( .IN1(n806), .IN2(rdata_1[14]), .IN3(n807), .IN4(rdata_0[14]), 
        .IN5(n1009), .Q(n1008) );
  AO22X1 U788 ( .IN1(n809), .IN2(rdata_2[14]), .IN3(n720), .IN4(rdata_7[14]), 
        .Q(n1009) );
  AO221X1 U789 ( .IN1(n810), .IN2(rdata_4[14]), .IN3(n811), .IN4(rdata_3[14]), 
        .IN5(n1010), .Q(n1007) );
  AO22X1 U790 ( .IN1(n813), .IN2(rdata_5[14]), .IN3(n814), .IN4(rdata_6[14]), 
        .Q(n1010) );
  NOR2X0 U791 ( .IN1(n713), .IN2(n760), .QN(N299) );
  NOR2X0 U792 ( .IN1(n713), .IN2(n761), .QN(N298) );
  NOR2X0 U793 ( .IN1(n713), .IN2(n762), .QN(N297) );
  NOR2X0 U794 ( .IN1(n713), .IN2(n763), .QN(N296) );
  NOR2X0 U795 ( .IN1(n713), .IN2(n764), .QN(N295) );
  NOR2X0 U796 ( .IN1(n713), .IN2(n765), .QN(N294) );
  NOR2X0 U797 ( .IN1(n713), .IN2(n766), .QN(N293) );
  NOR2X0 U798 ( .IN1(n713), .IN2(n767), .QN(N292) );
  NOR2X0 U799 ( .IN1(n713), .IN2(n768), .QN(N291) );
  NOR2X0 U800 ( .IN1(n713), .IN2(n769), .QN(N290) );
  OR2X1 U801 ( .IN1(n1011), .IN2(n1012), .Q(N29) );
  AO221X1 U802 ( .IN1(n806), .IN2(rdata_1[13]), .IN3(n807), .IN4(rdata_0[13]), 
        .IN5(n1013), .Q(n1012) );
  AO22X1 U803 ( .IN1(n809), .IN2(rdata_2[13]), .IN3(n720), .IN4(rdata_7[13]), 
        .Q(n1013) );
  AO221X1 U804 ( .IN1(n810), .IN2(rdata_4[13]), .IN3(n811), .IN4(rdata_3[13]), 
        .IN5(n1014), .Q(n1011) );
  AO22X1 U805 ( .IN1(n813), .IN2(rdata_5[13]), .IN3(n814), .IN4(rdata_6[13]), 
        .Q(n1014) );
  NOR2X0 U806 ( .IN1(n713), .IN2(n770), .QN(N289) );
  NOR2X0 U807 ( .IN1(n713), .IN2(n771), .QN(N288) );
  NOR2X0 U808 ( .IN1(n713), .IN2(n772), .QN(N287) );
  NOR2X0 U809 ( .IN1(n713), .IN2(n773), .QN(N286) );
  NOR2X0 U810 ( .IN1(n713), .IN2(n774), .QN(N285) );
  NOR2X0 U811 ( .IN1(n713), .IN2(n775), .QN(N284) );
  NOR2X0 U812 ( .IN1(n713), .IN2(n776), .QN(N283) );
  NOR2X0 U813 ( .IN1(n713), .IN2(n777), .QN(N282) );
  NOR2X0 U814 ( .IN1(n713), .IN2(n778), .QN(N281) );
  NOR2X0 U815 ( .IN1(n713), .IN2(n779), .QN(N280) );
  OR2X1 U816 ( .IN1(n1015), .IN2(n1016), .Q(N28) );
  AO221X1 U817 ( .IN1(n806), .IN2(rdata_1[12]), .IN3(n807), .IN4(rdata_0[12]), 
        .IN5(n1017), .Q(n1016) );
  AO22X1 U818 ( .IN1(n809), .IN2(rdata_2[12]), .IN3(n720), .IN4(rdata_7[12]), 
        .Q(n1017) );
  AO221X1 U819 ( .IN1(n810), .IN2(rdata_4[12]), .IN3(n811), .IN4(rdata_3[12]), 
        .IN5(n1018), .Q(n1015) );
  AO22X1 U820 ( .IN1(n813), .IN2(rdata_5[12]), .IN3(n814), .IN4(rdata_6[12]), 
        .Q(n1018) );
  NOR2X0 U821 ( .IN1(n713), .IN2(n780), .QN(N279) );
  NOR2X0 U822 ( .IN1(n713), .IN2(n781), .QN(N278) );
  NOR2X0 U823 ( .IN1(n713), .IN2(n782), .QN(N277) );
  NOR2X0 U824 ( .IN1(n713), .IN2(n783), .QN(N276) );
  NOR2X0 U825 ( .IN1(n713), .IN2(n784), .QN(N275) );
  NOR2X0 U826 ( .IN1(n713), .IN2(n785), .QN(N274) );
  NOR2X0 U827 ( .IN1(n713), .IN2(n786), .QN(N273) );
  NOR2X0 U828 ( .IN1(n803), .IN2(n723), .QN(N272) );
  NOR2X0 U829 ( .IN1(n803), .IN2(n724), .QN(N271) );
  NOR2X0 U830 ( .IN1(n803), .IN2(n725), .QN(N270) );
  OR2X1 U831 ( .IN1(n1019), .IN2(n1020), .Q(N27) );
  AO221X1 U832 ( .IN1(n806), .IN2(rdata_1[11]), .IN3(n807), .IN4(rdata_0[11]), 
        .IN5(n1021), .Q(n1020) );
  AO22X1 U833 ( .IN1(n809), .IN2(rdata_2[11]), .IN3(n720), .IN4(rdata_7[11]), 
        .Q(n1021) );
  AO221X1 U834 ( .IN1(n810), .IN2(rdata_4[11]), .IN3(n811), .IN4(rdata_3[11]), 
        .IN5(n1022), .Q(n1019) );
  AO22X1 U835 ( .IN1(n813), .IN2(rdata_5[11]), .IN3(n814), .IN4(rdata_6[11]), 
        .Q(n1022) );
  NOR2X0 U836 ( .IN1(n803), .IN2(n726), .QN(N269) );
  NOR2X0 U837 ( .IN1(n803), .IN2(n727), .QN(N268) );
  NOR2X0 U838 ( .IN1(n803), .IN2(n728), .QN(N267) );
  NOR2X0 U839 ( .IN1(n803), .IN2(n729), .QN(N266) );
  NOR2X0 U840 ( .IN1(n803), .IN2(n730), .QN(N265) );
  NOR2X0 U841 ( .IN1(n803), .IN2(n731), .QN(N264) );
  NOR2X0 U842 ( .IN1(n803), .IN2(n732), .QN(N263) );
  NOR2X0 U843 ( .IN1(n803), .IN2(n733), .QN(N262) );
  NOR2X0 U844 ( .IN1(n803), .IN2(n734), .QN(N261) );
  NOR2X0 U845 ( .IN1(n803), .IN2(n735), .QN(N260) );
  OR2X1 U846 ( .IN1(n1023), .IN2(n1024), .Q(N26) );
  AO221X1 U847 ( .IN1(n806), .IN2(rdata_1[10]), .IN3(n807), .IN4(rdata_0[10]), 
        .IN5(n1025), .Q(n1024) );
  AO22X1 U848 ( .IN1(n809), .IN2(rdata_2[10]), .IN3(n720), .IN4(rdata_7[10]), 
        .Q(n1025) );
  AO221X1 U849 ( .IN1(n810), .IN2(rdata_4[10]), .IN3(n811), .IN4(rdata_3[10]), 
        .IN5(n1026), .Q(n1023) );
  AO22X1 U850 ( .IN1(n813), .IN2(rdata_5[10]), .IN3(n814), .IN4(rdata_6[10]), 
        .Q(n1026) );
  NOR2X0 U851 ( .IN1(n803), .IN2(n736), .QN(N259) );
  NOR2X0 U852 ( .IN1(n803), .IN2(n737), .QN(N258) );
  NOR2X0 U853 ( .IN1(n803), .IN2(n738), .QN(N257) );
  NOR2X0 U854 ( .IN1(n803), .IN2(n739), .QN(N256) );
  NOR2X0 U855 ( .IN1(n803), .IN2(n740), .QN(N255) );
  NOR2X0 U856 ( .IN1(n803), .IN2(n741), .QN(N254) );
  NOR2X0 U857 ( .IN1(n803), .IN2(n742), .QN(N253) );
  NOR2X0 U858 ( .IN1(n803), .IN2(n743), .QN(N252) );
  NOR2X0 U859 ( .IN1(n803), .IN2(n744), .QN(N251) );
  NOR2X0 U860 ( .IN1(n803), .IN2(n745), .QN(N250) );
  OR2X1 U861 ( .IN1(n1027), .IN2(n1028), .Q(N25) );
  AO221X1 U862 ( .IN1(n806), .IN2(rdata_1[9]), .IN3(n807), .IN4(rdata_0[9]), 
        .IN5(n1029), .Q(n1028) );
  AO22X1 U863 ( .IN1(n809), .IN2(rdata_2[9]), .IN3(n720), .IN4(rdata_7[9]), 
        .Q(n1029) );
  AO221X1 U864 ( .IN1(n810), .IN2(rdata_4[9]), .IN3(n811), .IN4(rdata_3[9]), 
        .IN5(n1030), .Q(n1027) );
  AO22X1 U865 ( .IN1(n813), .IN2(rdata_5[9]), .IN3(n814), .IN4(rdata_6[9]), 
        .Q(n1030) );
  NOR2X0 U866 ( .IN1(n803), .IN2(n746), .QN(N249) );
  NOR2X0 U867 ( .IN1(n803), .IN2(n747), .QN(N248) );
  NOR2X0 U868 ( .IN1(n803), .IN2(n748), .QN(N247) );
  NOR2X0 U869 ( .IN1(n803), .IN2(n749), .QN(N246) );
  NOR2X0 U870 ( .IN1(n803), .IN2(n750), .QN(N245) );
  NOR2X0 U871 ( .IN1(n803), .IN2(n751), .QN(N244) );
  NOR2X0 U872 ( .IN1(n803), .IN2(n752), .QN(N243) );
  NOR2X0 U873 ( .IN1(n803), .IN2(n753), .QN(N242) );
  NOR2X0 U874 ( .IN1(n803), .IN2(n754), .QN(N241) );
  NOR2X0 U875 ( .IN1(n803), .IN2(n755), .QN(N240) );
  OR2X1 U876 ( .IN1(n1031), .IN2(n1032), .Q(N24) );
  AO221X1 U877 ( .IN1(n806), .IN2(rdata_1[8]), .IN3(n807), .IN4(rdata_0[8]), 
        .IN5(n1033), .Q(n1032) );
  AO22X1 U878 ( .IN1(n809), .IN2(rdata_2[8]), .IN3(n720), .IN4(rdata_7[8]), 
        .Q(n1033) );
  AO221X1 U879 ( .IN1(n810), .IN2(rdata_4[8]), .IN3(n811), .IN4(rdata_3[8]), 
        .IN5(n1034), .Q(n1031) );
  AO22X1 U880 ( .IN1(n813), .IN2(rdata_5[8]), .IN3(n814), .IN4(rdata_6[8]), 
        .Q(n1034) );
  NOR2X0 U881 ( .IN1(n803), .IN2(n756), .QN(N239) );
  NOR2X0 U882 ( .IN1(n803), .IN2(n757), .QN(N238) );
  NOR2X0 U883 ( .IN1(n803), .IN2(n758), .QN(N237) );
  NOR2X0 U884 ( .IN1(n803), .IN2(n759), .QN(N236) );
  NOR2X0 U885 ( .IN1(n803), .IN2(n760), .QN(N235) );
  NOR2X0 U886 ( .IN1(n803), .IN2(n761), .QN(N234) );
  NOR2X0 U887 ( .IN1(n803), .IN2(n762), .QN(N233) );
  NOR2X0 U888 ( .IN1(n803), .IN2(n763), .QN(N232) );
  NOR2X0 U889 ( .IN1(n803), .IN2(n764), .QN(N231) );
  NOR2X0 U890 ( .IN1(n803), .IN2(n765), .QN(N230) );
  OR2X1 U891 ( .IN1(n1035), .IN2(n1036), .Q(N23) );
  AO221X1 U892 ( .IN1(n806), .IN2(rdata_1[7]), .IN3(n807), .IN4(rdata_0[7]), 
        .IN5(n1037), .Q(n1036) );
  AO22X1 U893 ( .IN1(n809), .IN2(rdata_2[7]), .IN3(n720), .IN4(rdata_7[7]), 
        .Q(n1037) );
  AO221X1 U894 ( .IN1(n810), .IN2(rdata_4[7]), .IN3(n811), .IN4(rdata_3[7]), 
        .IN5(n1038), .Q(n1035) );
  AO22X1 U895 ( .IN1(n813), .IN2(rdata_5[7]), .IN3(n814), .IN4(rdata_6[7]), 
        .Q(n1038) );
  NOR2X0 U896 ( .IN1(n803), .IN2(n766), .QN(N229) );
  NOR2X0 U897 ( .IN1(n803), .IN2(n767), .QN(N228) );
  NOR2X0 U898 ( .IN1(n803), .IN2(n768), .QN(N227) );
  NOR2X0 U899 ( .IN1(n803), .IN2(n769), .QN(N226) );
  NOR2X0 U900 ( .IN1(n803), .IN2(n770), .QN(N225) );
  NOR2X0 U901 ( .IN1(n803), .IN2(n771), .QN(N224) );
  NOR2X0 U902 ( .IN1(n803), .IN2(n772), .QN(N223) );
  NOR2X0 U903 ( .IN1(n803), .IN2(n773), .QN(N222) );
  NOR2X0 U904 ( .IN1(n803), .IN2(n774), .QN(N221) );
  NOR2X0 U905 ( .IN1(n803), .IN2(n775), .QN(N220) );
  OR2X1 U906 ( .IN1(n1039), .IN2(n1040), .Q(N22) );
  AO221X1 U907 ( .IN1(n806), .IN2(rdata_1[6]), .IN3(n807), .IN4(rdata_0[6]), 
        .IN5(n1041), .Q(n1040) );
  AO22X1 U908 ( .IN1(n809), .IN2(rdata_2[6]), .IN3(n720), .IN4(rdata_7[6]), 
        .Q(n1041) );
  AO221X1 U909 ( .IN1(n810), .IN2(rdata_4[6]), .IN3(n811), .IN4(rdata_3[6]), 
        .IN5(n1042), .Q(n1039) );
  AO22X1 U910 ( .IN1(n813), .IN2(rdata_5[6]), .IN3(n814), .IN4(rdata_6[6]), 
        .Q(n1042) );
  NOR2X0 U911 ( .IN1(n803), .IN2(n776), .QN(N219) );
  NOR2X0 U912 ( .IN1(n803), .IN2(n777), .QN(N218) );
  NOR2X0 U913 ( .IN1(n803), .IN2(n778), .QN(N217) );
  NOR2X0 U914 ( .IN1(n803), .IN2(n779), .QN(N216) );
  NOR2X0 U915 ( .IN1(n803), .IN2(n780), .QN(N215) );
  NOR2X0 U916 ( .IN1(n803), .IN2(n781), .QN(N214) );
  NOR2X0 U917 ( .IN1(n803), .IN2(n782), .QN(N213) );
  NOR2X0 U918 ( .IN1(n803), .IN2(n783), .QN(N212) );
  NOR2X0 U919 ( .IN1(n803), .IN2(n784), .QN(N211) );
  NOR2X0 U920 ( .IN1(n803), .IN2(n785), .QN(N210) );
  OR2X1 U921 ( .IN1(n1043), .IN2(n1044), .Q(N21) );
  AO221X1 U922 ( .IN1(n806), .IN2(rdata_1[5]), .IN3(n807), .IN4(rdata_0[5]), 
        .IN5(n1045), .Q(n1044) );
  AO22X1 U923 ( .IN1(n809), .IN2(rdata_2[5]), .IN3(n720), .IN4(rdata_7[5]), 
        .Q(n1045) );
  AO221X1 U924 ( .IN1(n810), .IN2(rdata_4[5]), .IN3(n811), .IN4(rdata_3[5]), 
        .IN5(n1046), .Q(n1043) );
  AO22X1 U925 ( .IN1(n813), .IN2(rdata_5[5]), .IN3(n814), .IN4(rdata_6[5]), 
        .Q(n1046) );
  NOR2X0 U926 ( .IN1(n803), .IN2(n786), .QN(N209) );
  NOR2X0 U927 ( .IN1(n718), .IN2(n787), .QN(N208) );
  NOR2X0 U928 ( .IN1(n718), .IN2(n788), .QN(N207) );
  NOR2X0 U929 ( .IN1(n718), .IN2(n789), .QN(N206) );
  NOR2X0 U930 ( .IN1(n718), .IN2(n790), .QN(N205) );
  NOR2X0 U931 ( .IN1(n718), .IN2(n791), .QN(N204) );
  NOR2X0 U932 ( .IN1(n718), .IN2(n792), .QN(N203) );
  NOR2X0 U933 ( .IN1(n718), .IN2(n793), .QN(N202) );
  NOR2X0 U934 ( .IN1(n718), .IN2(n794), .QN(N201) );
  NOR2X0 U935 ( .IN1(n718), .IN2(n795), .QN(N200) );
  OR2X1 U936 ( .IN1(n1047), .IN2(n1048), .Q(N20) );
  AO221X1 U937 ( .IN1(n806), .IN2(rdata_1[4]), .IN3(n807), .IN4(rdata_0[4]), 
        .IN5(n1049), .Q(n1048) );
  AO22X1 U938 ( .IN1(n809), .IN2(rdata_2[4]), .IN3(n720), .IN4(rdata_7[4]), 
        .Q(n1049) );
  AO221X1 U939 ( .IN1(n810), .IN2(rdata_4[4]), .IN3(n811), .IN4(rdata_3[4]), 
        .IN5(n1050), .Q(n1047) );
  AO22X1 U940 ( .IN1(n813), .IN2(rdata_5[4]), .IN3(n814), .IN4(rdata_6[4]), 
        .Q(n1050) );
  NOR2X0 U941 ( .IN1(n718), .IN2(n796), .QN(N199) );
  NOR2X0 U942 ( .IN1(n718), .IN2(n797), .QN(N198) );
  NOR2X0 U943 ( .IN1(n718), .IN2(n798), .QN(N197) );
  NOR2X0 U944 ( .IN1(n718), .IN2(n799), .QN(N196) );
  NOR2X0 U945 ( .IN1(n718), .IN2(n800), .QN(N195) );
  NOR2X0 U946 ( .IN1(n718), .IN2(n801), .QN(N194) );
  NOR2X0 U947 ( .IN1(n718), .IN2(n802), .QN(N193) );
  NOR2X0 U948 ( .IN1(n719), .IN2(n787), .QN(N192) );
  NOR2X0 U949 ( .IN1(n719), .IN2(n788), .QN(N191) );
  NOR2X0 U950 ( .IN1(n719), .IN2(n789), .QN(N190) );
  OR2X1 U951 ( .IN1(n1051), .IN2(n1052), .Q(N19) );
  AO221X1 U952 ( .IN1(n806), .IN2(rdata_1[3]), .IN3(n807), .IN4(rdata_0[3]), 
        .IN5(n1053), .Q(n1052) );
  AO22X1 U953 ( .IN1(n809), .IN2(rdata_2[3]), .IN3(n720), .IN4(rdata_7[3]), 
        .Q(n1053) );
  AO221X1 U954 ( .IN1(n810), .IN2(rdata_4[3]), .IN3(n811), .IN4(rdata_3[3]), 
        .IN5(n1054), .Q(n1051) );
  AO22X1 U955 ( .IN1(n813), .IN2(rdata_5[3]), .IN3(n814), .IN4(rdata_6[3]), 
        .Q(n1054) );
  NOR2X0 U956 ( .IN1(n719), .IN2(n790), .QN(N189) );
  NOR2X0 U957 ( .IN1(n719), .IN2(n791), .QN(N188) );
  NOR2X0 U958 ( .IN1(n719), .IN2(n792), .QN(N187) );
  NOR2X0 U959 ( .IN1(n719), .IN2(n793), .QN(N186) );
  NOR2X0 U960 ( .IN1(n719), .IN2(n794), .QN(N185) );
  NOR2X0 U961 ( .IN1(n719), .IN2(n795), .QN(N184) );
  NOR2X0 U962 ( .IN1(n719), .IN2(n796), .QN(N183) );
  NOR2X0 U963 ( .IN1(n719), .IN2(n797), .QN(N182) );
  NOR2X0 U964 ( .IN1(n719), .IN2(n798), .QN(N181) );
  NOR2X0 U965 ( .IN1(n719), .IN2(n799), .QN(N180) );
  OR2X1 U966 ( .IN1(n1055), .IN2(n1056), .Q(N18) );
  AO221X1 U967 ( .IN1(n806), .IN2(rdata_1[2]), .IN3(n807), .IN4(rdata_0[2]), 
        .IN5(n1057), .Q(n1056) );
  AO22X1 U968 ( .IN1(n809), .IN2(rdata_2[2]), .IN3(n720), .IN4(rdata_7[2]), 
        .Q(n1057) );
  AO221X1 U969 ( .IN1(n810), .IN2(rdata_4[2]), .IN3(n811), .IN4(rdata_3[2]), 
        .IN5(n1058), .Q(n1055) );
  AO22X1 U970 ( .IN1(n813), .IN2(rdata_5[2]), .IN3(n814), .IN4(rdata_6[2]), 
        .Q(n1058) );
  NOR2X0 U971 ( .IN1(n719), .IN2(n800), .QN(N179) );
  NOR2X0 U972 ( .IN1(n719), .IN2(n801), .QN(N178) );
  NOR2X0 U973 ( .IN1(n719), .IN2(n802), .QN(N177) );
  NOR2X0 U974 ( .IN1(n717), .IN2(n787), .QN(N176) );
  NOR2X0 U975 ( .IN1(n717), .IN2(n788), .QN(N175) );
  NOR2X0 U976 ( .IN1(n717), .IN2(n789), .QN(N174) );
  NOR2X0 U977 ( .IN1(n717), .IN2(n790), .QN(N173) );
  NOR2X0 U978 ( .IN1(n717), .IN2(n791), .QN(N172) );
  NOR2X0 U979 ( .IN1(n717), .IN2(n792), .QN(N171) );
  NOR2X0 U980 ( .IN1(n717), .IN2(n793), .QN(N170) );
  OR2X1 U981 ( .IN1(n1059), .IN2(n1060), .Q(N17) );
  AO221X1 U982 ( .IN1(n806), .IN2(rdata_1[1]), .IN3(n807), .IN4(rdata_0[1]), 
        .IN5(n1061), .Q(n1060) );
  AO22X1 U983 ( .IN1(n809), .IN2(rdata_2[1]), .IN3(n720), .IN4(rdata_7[1]), 
        .Q(n1061) );
  AO221X1 U984 ( .IN1(n810), .IN2(rdata_4[1]), .IN3(n811), .IN4(rdata_3[1]), 
        .IN5(n1062), .Q(n1059) );
  AO22X1 U985 ( .IN1(n813), .IN2(rdata_5[1]), .IN3(n814), .IN4(rdata_6[1]), 
        .Q(n1062) );
  NOR2X0 U986 ( .IN1(n717), .IN2(n794), .QN(N169) );
  NOR2X0 U987 ( .IN1(n717), .IN2(n795), .QN(N168) );
  NOR2X0 U988 ( .IN1(n717), .IN2(n796), .QN(N167) );
  NOR2X0 U989 ( .IN1(n717), .IN2(n797), .QN(N166) );
  NOR2X0 U990 ( .IN1(n717), .IN2(n798), .QN(N165) );
  NOR2X0 U991 ( .IN1(n717), .IN2(n799), .QN(N164) );
  NOR2X0 U992 ( .IN1(n717), .IN2(n800), .QN(N163) );
  NOR2X0 U993 ( .IN1(n717), .IN2(n801), .QN(N162) );
  NOR2X0 U994 ( .IN1(n717), .IN2(n802), .QN(N161) );
  NOR2X0 U995 ( .IN1(n715), .IN2(n787), .QN(N160) );
  OR2X1 U996 ( .IN1(n1063), .IN2(n1064), .Q(N16) );
  AO221X1 U997 ( .IN1(n806), .IN2(rdata_1[0]), .IN3(n807), .IN4(rdata_0[0]), 
        .IN5(n1065), .Q(n1064) );
  AO22X1 U998 ( .IN1(n809), .IN2(rdata_2[0]), .IN3(n720), .IN4(rdata_7[0]), 
        .Q(n1065) );
  AO221X1 U1004 ( .IN1(n810), .IN2(rdata_4[0]), .IN3(n811), .IN4(rdata_3[0]), 
        .IN5(n1067), .Q(n1063) );
  AO22X1 U1005 ( .IN1(n813), .IN2(rdata_5[0]), .IN3(n814), .IN4(rdata_6[0]), 
        .Q(n1067) );
  NOR2X0 U1006 ( .IN1(n715), .IN2(n788), .QN(N159) );
  NOR2X0 U1007 ( .IN1(n715), .IN2(n789), .QN(N158) );
  NOR2X0 U1008 ( .IN1(n715), .IN2(n790), .QN(N157) );
  NOR2X0 U1009 ( .IN1(n715), .IN2(n791), .QN(N156) );
  NOR2X0 U1010 ( .IN1(n715), .IN2(n792), .QN(N155) );
  NOR2X0 U1011 ( .IN1(n715), .IN2(n793), .QN(N154) );
  NOR2X0 U1012 ( .IN1(n715), .IN2(n794), .QN(N153) );
  NOR2X0 U1013 ( .IN1(n715), .IN2(n795), .QN(N152) );
  NOR2X0 U1014 ( .IN1(n715), .IN2(n796), .QN(N151) );
  NOR2X0 U1015 ( .IN1(n715), .IN2(n797), .QN(N150) );
  NOR2X0 U1016 ( .IN1(n715), .IN2(n798), .QN(N149) );
  NOR2X0 U1017 ( .IN1(n715), .IN2(n799), .QN(N148) );
  NOR2X0 U1018 ( .IN1(n715), .IN2(n800), .QN(N147) );
  NOR2X0 U1019 ( .IN1(n715), .IN2(n801), .QN(N146) );
  NOR2X0 U1020 ( .IN1(n715), .IN2(n802), .QN(N145) );
  NOR2X0 U1023 ( .IN1(n716), .IN2(n787), .QN(N144) );
  NOR2X0 U1024 ( .IN1(n716), .IN2(n788), .QN(N143) );
  NOR2X0 U1025 ( .IN1(n716), .IN2(n789), .QN(N142) );
  NOR2X0 U1026 ( .IN1(n716), .IN2(n790), .QN(N141) );
  NOR2X0 U1027 ( .IN1(n716), .IN2(n791), .QN(N140) );
  NOR2X0 U1028 ( .IN1(n716), .IN2(n792), .QN(N139) );
  NOR2X0 U1029 ( .IN1(n716), .IN2(n793), .QN(N138) );
  NOR2X0 U1030 ( .IN1(n716), .IN2(n794), .QN(N137) );
  NOR2X0 U1031 ( .IN1(n716), .IN2(n795), .QN(N136) );
  NOR2X0 U1032 ( .IN1(n716), .IN2(n796), .QN(N135) );
  NOR2X0 U1033 ( .IN1(n716), .IN2(n797), .QN(N134) );
  NOR2X0 U1034 ( .IN1(n716), .IN2(n798), .QN(N133) );
  NOR2X0 U1035 ( .IN1(n716), .IN2(n799), .QN(N132) );
  NOR2X0 U1036 ( .IN1(n716), .IN2(n800), .QN(N131) );
  NOR2X0 U1037 ( .IN1(n716), .IN2(n801), .QN(N130) );
  NOR2X0 U1038 ( .IN1(n716), .IN2(n802), .QN(N129) );
  NOR2X0 U1041 ( .IN1(n714), .IN2(n787), .QN(N128) );
  NOR2X0 U1042 ( .IN1(n714), .IN2(n788), .QN(N127) );
  NOR2X0 U1043 ( .IN1(n714), .IN2(n789), .QN(N126) );
  NOR2X0 U1044 ( .IN1(n714), .IN2(n790), .QN(N125) );
  NOR2X0 U1045 ( .IN1(n714), .IN2(n791), .QN(N124) );
  NOR2X0 U1046 ( .IN1(n714), .IN2(n792), .QN(N123) );
  NOR2X0 U1047 ( .IN1(n714), .IN2(n793), .QN(N122) );
  NOR2X0 U1048 ( .IN1(n714), .IN2(n794), .QN(N121) );
  NOR2X0 U1049 ( .IN1(n714), .IN2(n795), .QN(N120) );
  NOR2X0 U1050 ( .IN1(n714), .IN2(n796), .QN(N119) );
  NOR2X0 U1051 ( .IN1(n714), .IN2(n797), .QN(N118) );
  NOR2X0 U1052 ( .IN1(n714), .IN2(n798), .QN(N117) );
  NOR2X0 U1053 ( .IN1(n714), .IN2(n799), .QN(N116) );
  NOR2X0 U1054 ( .IN1(n714), .IN2(n800), .QN(N115) );
  NOR2X0 U1055 ( .IN1(n714), .IN2(n801), .QN(N114) );
  NOR2X0 U1056 ( .IN1(n714), .IN2(n802), .QN(N113) );
  NOR2X0 U1059 ( .IN1(n713), .IN2(n787), .QN(N112) );
  NOR2X0 U1060 ( .IN1(n713), .IN2(n788), .QN(N111) );
  NOR2X0 U1061 ( .IN1(n713), .IN2(n789), .QN(N110) );
  NOR2X0 U1062 ( .IN1(n713), .IN2(n790), .QN(N109) );
  NOR2X0 U1063 ( .IN1(n713), .IN2(n791), .QN(N108) );
  NOR2X0 U1064 ( .IN1(n713), .IN2(n792), .QN(N107) );
  NOR2X0 U1065 ( .IN1(n713), .IN2(n793), .QN(N106) );
  NOR2X0 U1066 ( .IN1(n713), .IN2(n794), .QN(N105) );
  NOR2X0 U1067 ( .IN1(n713), .IN2(n795), .QN(N104) );
  NOR2X0 U1068 ( .IN1(n713), .IN2(n796), .QN(N103) );
  NOR2X0 U1069 ( .IN1(n713), .IN2(n797), .QN(N102) );
  NOR2X0 U1070 ( .IN1(n713), .IN2(n798), .QN(N101) );
  NOR2X0 U1071 ( .IN1(n713), .IN2(n799), .QN(N100) );
  INVX0 U67 ( .IN(wdata_mbist[9]), .QN(n777) );
  INVX0 U66 ( .IN(wdata_mbist[10]), .QN(n776) );
  INVX0 U69 ( .IN(wdata_mbist[7]), .QN(n779) );
  INVX0 U70 ( .IN(wdata_mbist[6]), .QN(n780) );
  INVX0 U75 ( .IN(wdata_mbist[1]), .QN(n785) );
  INVX0 U71 ( .IN(wdata_mbist[5]), .QN(n781) );
  INVX0 U72 ( .IN(wdata_mbist[4]), .QN(n782) );
  INVX0 U73 ( .IN(wdata_mbist[3]), .QN(n783) );
  INVX0 U74 ( .IN(wdata_mbist[2]), .QN(n784) );
  INVX0 U68 ( .IN(wdata_mbist[8]), .QN(n778) );
  INVX0 U65 ( .IN(wdata_mbist[11]), .QN(n775) );
  INVX0 U64 ( .IN(wdata_mbist[12]), .QN(n774) );
  INVX0 U63 ( .IN(wdata_mbist[13]), .QN(n773) );
  INVX0 U62 ( .IN(wdata_mbist[14]), .QN(n772) );
  INVX0 U61 ( .IN(wdata_mbist[15]), .QN(n771) );
  INVX0 U60 ( .IN(wdata_mbist[16]), .QN(n770) );
  INVX0 U59 ( .IN(wdata_mbist[17]), .QN(n769) );
  INVX0 U58 ( .IN(wdata_mbist[18]), .QN(n768) );
  INVX0 U57 ( .IN(wdata_mbist[19]), .QN(n767) );
  INVX0 U56 ( .IN(wdata_mbist[20]), .QN(n766) );
  INVX0 U54 ( .IN(wdata_mbist[22]), .QN(n764) );
  INVX0 U53 ( .IN(wdata_mbist[23]), .QN(n763) );
  INVX0 U52 ( .IN(wdata_mbist[24]), .QN(n762) );
  INVX0 U51 ( .IN(wdata_mbist[25]), .QN(n761) );
  INVX0 U50 ( .IN(wdata_mbist[26]), .QN(n760) );
  INVX0 U49 ( .IN(wdata_mbist[27]), .QN(n759) );
  INVX0 U48 ( .IN(wdata_mbist[28]), .QN(n758) );
  INVX0 U47 ( .IN(wdata_mbist[29]), .QN(n757) );
  INVX0 U46 ( .IN(wdata_mbist[30]), .QN(n756) );
  INVX0 U45 ( .IN(wdata_mbist[31]), .QN(n755) );
  INVX0 U44 ( .IN(wdata_mbist[32]), .QN(n754) );
  INVX0 U43 ( .IN(wdata_mbist[33]), .QN(n753) );
  INVX0 U42 ( .IN(wdata_mbist[34]), .QN(n752) );
  INVX0 U41 ( .IN(wdata_mbist[35]), .QN(n751) );
  INVX0 U40 ( .IN(wdata_mbist[36]), .QN(n750) );
  INVX0 U39 ( .IN(wdata_mbist[37]), .QN(n749) );
  INVX0 U38 ( .IN(wdata_mbist[38]), .QN(n748) );
  INVX0 U37 ( .IN(wdata_mbist[39]), .QN(n747) );
  INVX0 U36 ( .IN(wdata_mbist[40]), .QN(n746) );
  INVX0 U35 ( .IN(wdata_mbist[41]), .QN(n745) );
  INVX0 U34 ( .IN(wdata_mbist[42]), .QN(n744) );
  INVX0 U33 ( .IN(wdata_mbist[43]), .QN(n743) );
  INVX0 U32 ( .IN(wdata_mbist[44]), .QN(n742) );
  INVX0 U31 ( .IN(wdata_mbist[45]), .QN(n741) );
  INVX0 U30 ( .IN(wdata_mbist[46]), .QN(n740) );
  INVX0 U29 ( .IN(wdata_mbist[47]), .QN(n739) );
  INVX0 U28 ( .IN(wdata_mbist[48]), .QN(n738) );
  INVX0 U27 ( .IN(wdata_mbist[49]), .QN(n737) );
  INVX0 U26 ( .IN(wdata_mbist[50]), .QN(n736) );
  INVX0 U25 ( .IN(wdata_mbist[51]), .QN(n735) );
  INVX0 U24 ( .IN(wdata_mbist[52]), .QN(n734) );
  INVX0 U23 ( .IN(wdata_mbist[53]), .QN(n733) );
  INVX0 U22 ( .IN(wdata_mbist[54]), .QN(n732) );
  INVX0 U21 ( .IN(wdata_mbist[55]), .QN(n731) );
  INVX0 U20 ( .IN(wdata_mbist[56]), .QN(n730) );
  INVX0 U19 ( .IN(wdata_mbist[57]), .QN(n729) );
  INVX0 U18 ( .IN(wdata_mbist[58]), .QN(n728) );
  INVX0 U17 ( .IN(wdata_mbist[59]), .QN(n727) );
  INVX0 U55 ( .IN(wdata_mbist[21]), .QN(n765) );
  INVX0 U16 ( .IN(wdata_mbist[60]), .QN(n726) );
  INVX0 U76 ( .IN(wdata_mbist[0]), .QN(n786) );
  INVX0 U14 ( .IN(wdata_mbist[62]), .QN(n724) );
  INVX0 U13 ( .IN(wdata_mbist[63]), .QN(n723) );
  INVX0 U15 ( .IN(wdata_mbist[61]), .QN(n725) );
  INVX0 U11 ( .IN(memory_sel[0]), .QN(n721) );
  INVX0 U88 ( .IN(address_mbist[4]), .QN(n798) );
  INVX0 U87 ( .IN(address_mbist[5]), .QN(n797) );
  INVX0 U86 ( .IN(address_mbist[6]), .QN(n796) );
  INVX0 U85 ( .IN(address_mbist[7]), .QN(n795) );
  INVX0 U84 ( .IN(address_mbist[8]), .QN(n794) );
  INVX0 U83 ( .IN(address_mbist[9]), .QN(n793) );
  INVX0 U82 ( .IN(address_mbist[10]), .QN(n792) );
  INVX0 U12 ( .IN(write_read_mbist), .QN(n722) );
  INVX0 U81 ( .IN(address_mbist[11]), .QN(n791) );
  INVX0 U80 ( .IN(address_mbist[12]), .QN(n790) );
  INVX0 U79 ( .IN(address_mbist[13]), .QN(n789) );
  INVX0 U78 ( .IN(address_mbist[14]), .QN(n788) );
  INVX0 U77 ( .IN(address_mbist[15]), .QN(n787) );
  INVX0 U91 ( .IN(address_mbist[1]), .QN(n801) );
  INVX0 U90 ( .IN(address_mbist[2]), .QN(n800) );
  INVX0 U89 ( .IN(address_mbist[3]), .QN(n799) );
  INVX0 U92 ( .IN(address_mbist[0]), .QN(n802) );
  NOR3X0 U1003 ( .IN1(memory_sel[2]), .IN2(memory_sel[1]), .IN3(n721), .QN(
        n806) );
  NOR3X0 U1002 ( .IN1(memory_sel[0]), .IN2(memory_sel[2]), .IN3(memory_sel[1]), 
        .QN(n807) );
  NOR2X0 U1072 ( .IN1(memory_sel[0]), .IN2(n1071), .QN(n814) );
  NAND3X0 U999 ( .IN1(memory_sel[0]), .IN2(memory_sel[2]), .IN3(memory_sel[1]), 
        .QN(n803) );
  NOR2X0 U1039 ( .IN1(memory_sel[1]), .IN2(n1069), .QN(n810) );
  NOR2X0 U1021 ( .IN1(memory_sel[2]), .IN2(n1068), .QN(n811) );
  NOR2X0 U1000 ( .IN1(memory_sel[2]), .IN2(n1066), .QN(n809) );
  NOR2X0 U1057 ( .IN1(memory_sel[1]), .IN2(n1070), .QN(n813) );
  NAND2X0 U1073 ( .IN1(memory_sel[2]), .IN2(memory_sel[1]), .QN(n1071) );
  NAND2X0 U1058 ( .IN1(memory_sel[0]), .IN2(memory_sel[2]), .QN(n1070) );
  NAND2X0 U1022 ( .IN1(memory_sel[0]), .IN2(memory_sel[1]), .QN(n1068) );
  NAND2X0 U1040 ( .IN1(memory_sel[2]), .IN2(n721), .QN(n1069) );
  NAND2X0 U1001 ( .IN1(memory_sel[1]), .IN2(n721), .QN(n1066) );
  INVX0 U3 ( .IN(n814), .QN(n713) );
  INVX0 U4 ( .IN(n813), .QN(n714) );
  INVX0 U5 ( .IN(n809), .QN(n717) );
  INVX0 U6 ( .IN(n811), .QN(n715) );
  INVX0 U7 ( .IN(n807), .QN(n718) );
  INVX0 U8 ( .IN(n810), .QN(n716) );
  INVX0 U9 ( .IN(n806), .QN(n719) );
  INVX0 U10 ( .IN(n803), .QN(n720) );
endmodule


module vr ( clk, rst_n, test_mode, operation, error_exceed_ignore, 
        allowable_faulty, memory_sel, address_7, address_6, address_5, 
        address_4, address_3, address_2, address_1, address_0, write_read_7, 
        write_read_6, write_read_5, write_read_4, write_read_3, write_read_2, 
        write_read_1, write_read_0, memtype, wdata_7, wdata_6, wdata_5, 
        wdata_4, wdata_3, wdata_2, wdata_1, wdata_0, rdata_7, rdata_6, rdata_5, 
        rdata_4, rdata_3, rdata_2, rdata_1, rdata_0, error, force_terminate, 
        complete );
  input [2:0] operation;
  input [15:0] allowable_faulty;
  input [2:0] memory_sel;
  output [15:0] address_7;
  output [15:0] address_6;
  output [15:0] address_5;
  output [15:0] address_4;
  output [15:0] address_3;
  output [15:0] address_2;
  output [15:0] address_1;
  output [15:0] address_0;
  input [4:0] memtype;
  output [63:0] wdata_7;
  output [63:0] wdata_6;
  output [63:0] wdata_5;
  output [63:0] wdata_4;
  output [63:0] wdata_3;
  output [63:0] wdata_2;
  output [63:0] wdata_1;
  output [63:0] wdata_0;
  input [63:0] rdata_7;
  input [63:0] rdata_6;
  input [63:0] rdata_5;
  input [63:0] rdata_4;
  input [63:0] rdata_3;
  input [63:0] rdata_2;
  input [63:0] rdata_1;
  input [63:0] rdata_0;
  input clk, rst_n, test_mode, error_exceed_ignore;
  output write_read_7, write_read_6, write_read_5, write_read_4, write_read_3,
         write_read_2, write_read_1, write_read_0, error, force_terminate,
         complete;
  wire   anpsf_complete, apnpsf_en, write_read;
  wire   [15:0] address;
  wire   [63:0] wdata;
  wire   [63:0] rdata;

  controller controller_1 ( .clk(clk), .rst_n(rst_n), .test_mode(test_mode), 
        .operation({1'b0, 1'b0, 1'b0}), .apnpsf_complete(anpsf_complete), 
        .apnpsf_en(apnpsf_en), .complete(complete) );
  mbist_decoder mbist_decoder_1 ( .clk(clk), .rst_n(rst_n), .apnpsf_en(
        apnpsf_en), .error_exceed_ignore(error_exceed_ignore), 
        .allowable_faulty(allowable_faulty), .memtype(memtype), .address(
        address), .write_read(write_read), .wdata(wdata), .rdata(rdata), 
        .error(error), .force_terminate(force_terminate), .apnpsf_complete(
        anpsf_complete) );
  mbist_mux_demux mbist_mux_demux_1 ( .clk(clk), .rst_n(rst_n), .memory_sel(
        memory_sel), .write_read_mbist(write_read), .rdata_mbist(rdata), 
        .wdata_mbist(wdata), .address_mbist(address), .write_read_7(
        write_read_7), .write_read_6(write_read_6), .write_read_5(write_read_5), .write_read_4(write_read_4), .write_read_3(write_read_3), .write_read_2(
        write_read_2), .write_read_1(write_read_1), .write_read_0(write_read_0), .rdata_7(rdata_7), .rdata_6(rdata_6), .rdata_5(rdata_5), .rdata_4(rdata_4), 
        .rdata_3(rdata_3), .rdata_2(rdata_2), .rdata_1(rdata_1), .rdata_0(
        rdata_0), .wdata_7(wdata_7), .wdata_6(wdata_6), .wdata_5(wdata_5), 
        .wdata_4(wdata_4), .wdata_3(wdata_3), .wdata_2(wdata_2), .wdata_1(
        wdata_1), .wdata_0(wdata_0), .address_7(address_7), .address_6(
        address_6), .address_5(address_5), .address_4(address_4), .address_3(
        address_3), .address_2(address_2), .address_1(address_1), .address_0(
        address_0) );
endmodule

